name C7552.iscas
i 1(0)
i 5(1)
i 9(2)
i 12(3)
i 15(4)
i 18(5)
i 23(6)
i 26(7)
i 29(8)
i 32(9)
i 35(10)
i 38(11)
i 41(12)
i 44(13)
i 47(14)
i 50(15)
i 53(16)
i 54(17)
i 55(18)
i 56(19)
i 57(20)
i 58(21)
i 59(22)
i 60(23)
i 61(24)
i 62(25)
i 63(26)
i 64(27)
i 65(28)
i 66(29)
i 69(30)
i 70(31)
i 73(32)
i 74(33)
i 75(34)
i 76(35)
i 77(36)
i 78(37)
i 79(38)
i 80(39)
i 81(40)
i 82(41)
i 83(42)
i 84(43)
i 85(44)
i 86(45)
i 87(46)
i 88(47)
i 89(48)
i 94(49)
i 97(50)
i 100(51)
i 103(52)
i 106(53)
i 109(54)
i 110(55)
i 111(56)
i 112(57)
i 113(58)
i 114(59)
i 115(60)
i 118(61)
i 121(62)
i 124(63)
i 127(64)
i 130(65)
i 133(66)
i 134(67)
i 135(68)
i 138(69)
i 141(70)
i 144(71)
i 147(72)
i 150(73)
i 151(74)
i 152(75)
i 153(76)
i 154(77)
i 155(78)
i 156(79)
i 157(80)
i 158(81)
i 159(82)
i 160(83)
i 161(84)
i 162(85)
i 163(86)
i 164(87)
i 165(88)
i 166(89)
i 167(90)
i 168(91)
i 169(92)
i 170(93)
i 171(94)
i 172(95)
i 173(96)
i 174(97)
i 175(98)
i 176(99)
i 177(100)
i 178(101)
i 179(102)
i 180(103)
i 181(104)
i 182(105)
i 183(106)
i 184(107)
i 185(108)
i 186(109)
i 187(110)
i 188(111)
i 189(112)
i 190(113)
i 191(114)
i 192(115)
i 193(116)
i 194(117)
i 195(118)
i 196(119)
i 197(120)
i 198(121)
i 199(122)
i 200(123)
i 201(124)
i 202(125)
i 203(126)
i 204(127)
i 205(128)
i 206(129)
i 207(130)
i 208(131)
i 209(132)
i 210(133)
i 211(134)
i 212(135)
i 213(136)
i 214(137)
i 215(138)
i 216(139)
i 217(140)
i 218(141)
i 219(142)
i 220(143)
i 221(144)
i 222(145)
i 223(146)
i 224(147)
i 225(148)
i 226(149)
i 227(150)
i 228(151)
i 229(152)
i 230(153)
i 231(154)
i 232(155)
i 233(156)
i 234(157)
i 235(158)
i 236(159)
i 237(160)
i 238(161)
i 239(162)
i 240(163)
i IN-339(164)
i 1197(165)
i 1455(166)
i 1459(167)
i 1462(168)
i 1469(169)
i 1480(170)
i 1486(171)
i 1492(172)
i 1496(173)
i 2204(174)
i 2208(175)
i 2211(176)
i 2218(177)
i 2224(178)
i 2230(179)
i 2236(180)
i 2239(181)
i 2247(182)
i 2253(183)
i 2256(184)
i 3698(185)
i 3701(186)
i 3705(187)
i 3711(188)
i 3717(189)
i 3723(190)
i 3729(191)
i 3737(192)
i 3743(193)
i 3749(194)
i 4393(195)
i 4394(196)
i 4400(197)
i 4405(198)
i 4410(199)
i 4415(200)
i 4420(201)
i 4427(202)
i 4432(203)
i 4437(204)
i 4526(205)
i 4528(206)

o 339(164)
o 2(313)
o 3(312)
o 450(288)
o 448(284)
o 444(282)
o 442(280)
o 440(277)
o 438(274)
o 496(271)
o 494(267)
o 492(265)
o 490(263)
o 488(260)
o 486(258)
o 484(256)
o 482(253)
o 480(250)
o 560(248)
o 542(246)
o 558(244)
o 556(242)
o 554(240)
o 552(238)
o 550(236)
o 548(234)
o 546(232)
o 544(230)
o 540(227)
o 538(224)
o 536(222)
o 534(220)
o 532(218)
o 530(216)
o 528(214)
o 526(212)
o 524(210)
o 279(304)
o 436(286)
o 478(269)
o 522(226)
o 402(395)
o 404(390)
o 406(388)
o 408(385)
o 410(387)
o 432(428)
o 446(393)
o 284(384)
o 286(419)
o 289(383)
o 292(392)
o 341(420)
o 281(547)
o 453(596)
o 278(536)
o 373(2994)
o 246(3110)
o 258(3122)
o 264(3121)
o 270(3109)
o 388(3093)
o 391(3094)
o 394(3095)
o 397(3097)
o 376(3206)
o 379(3207)
o 382(3148)
o 385(3151)
o 412(3369)
o 414(3338)
o 416(3368)
o 249(3418)
o 295(3352)
o 324(3363)
o 252(3450)
o 276(3401)
o 310(3393)
o 313(3396)
o 316(3397)
o 319(3398)
o 327(3408)
o 330(3411)
o 333(3416)
o 336(3412)
o 418(3449)
o 273(3402)
o 298(3387)
o 301(3388)
o 304(3390)
o 307(3389)
o 344(3382)
o 422(3451)
o 469(3452)
o 419(3444)
o 471(3445)
o 359(3426)
o 362(3429)
o 365(3430)
o 368(3431)
o 347(3420)
o 350(3421)
o 353(3425)
o 356(3424)
o 321(3715)
o 338(3716)
o 370(3718)
o 399(3717)

g1 not 15(4) ; 279(304)
g2 or 401(310)* 400(297)* ; 402(395)
g3 not 2857(293) ; 404(390)
g4 not 4514(292) ; 406(388)
g5 not 4442(290) ; 408(385)
g6 not 1501(291) ; 410(387)
g7 or 574(308)* 1197(165)* ; 284(384)
g8 not 1205(305) ; 286(419)
g9 or 574(308)* 1197(165)* ; 289(383)
g10 or 575(309)* 1184(294)* ; 292(392)
g11 not 1205(305) ; 341(420)
g12 not 280(391) ; 281(547)
g13 and 453(596) 163(86) ; 278(536)
g14 or 372(2890)* 371(2754)* ; 373(2994)
g15 or 245(2897) 244(3033) 243(3032) 242(2955) 241(2837) ; 246(3110)
g16 or 257(2860) 256(2991) 255(2990) 254(2888) 3259(2874) ; 258(3122)
g17 or 263(2858) 262(2993) 261(2992) 260(2889) 3259(2874) ; 264(3121)
g18 or 269(2896) 268(3028) 267(3027) 266(2956) 265(2835) ; 270(3109)
g19 or 387(2931)* 386(3020)* ; 388(3093)
g20 or 390(2934)* 389(3021)* ; 391(3094)
g21 or 393(2937)* 392(3022)* ; 394(3095)
g22 or 396(2941)* 395(3023)* ; 397(3097)
g23 or 375(3090) 374(3152) ; 376(3206)
g24 or 378(3091) 377(3153) ; 379(3207)
g25 or 381(3092) 380(3086) ; 382(3148)
g26 or 384(3016) 383(3089) ; 385(3151)
g27 not 4443(3309) ; 412(3369)
g28 not 4524(3265) ; 414(3338)
g29 not 2868(3308) ; 416(3368)
g30 or 248(3306) 247(3310) ; 249(3418)
g31 or 294(3223)* 293(3285)* ; 295(3352)
g32 or 323(3238)* 322(3302)* ; 324(3363)
g33 or 251(3365) 250(3417) ; 252(3450)
g34 or 275(3286) 274(3353) ; 276(3401)
g35 or 309(3275)* 308(3346)* ; 310(3393)
g36 or 312(3279)* 311(3349)* ; 313(3396)
g37 or 315(3281)* 314(3350)* ; 316(3397)
g38 or 318(3283)* 317(3351)* ; 319(3398)
g39 or 326(3294)* 325(3358)* ; 327(3408)
g40 or 329(3298)* 328(3361)* ; 330(3411)
g41 or 332(3304)* 331(3364)* ; 333(3416)
g42 or 335(3300)* 334(3362)* ; 336(3412)
g43 not 417(3415) ; 418(3449)
g44 or 272(3287) 271(3354) ; 273(3402)
g45 or 297(3266) 296(3340) ; 298(3387)
g46 or 300(3267) 299(3341) ; 301(3388)
g47 or 303(3271) 302(3342) ; 304(3390)
g48 or 306(3270) 305(3343) ; 307(3389)
g49 or 343(3258)* 342(3330)* ; 344(3382)
g50 or 358(3320)* 357(3376)* ; 359(3426)
g51 or 361(3324)* 360(3379)* ; 362(3429)
g52 or 364(3326)* 363(3380)* ; 365(3430)
g53 or 367(3328)* 366(3381)* ; 368(3431)
g54 or 346(3311) 345(3370) ; 347(3420)
g55 or 349(3314) 348(3371) ; 350(3421)
g56 or 352(3318) 351(3372) ; 353(3425)
g57 or 355(3317) 354(3375) ; 356(3424)
g58 not 320(3711) ; 321(3715)
g59 not 337(3712) ; 338(3716)
g60 not 369(3714) ; 370(3718)
g61 not 398(3713) ; 399(3717)
g62 and 4526(205) ; 4833(207)
g63 and 4526(205) ; 2828(208)
g64 not 4437(204) ; 4439(209)
g65 not 4432(203) ; 4434(211)
g66 not 4427(202) ; 4429(213)
g67 not 4420(201) ; 4422(215)
g68 not 4415(200) ; 4417(217)
g69 not 4410(199) ; 4412(219)
g70 not 4405(198) ; 4407(221)
g71 not 4400(197) ; 4402(223)
g72 not 4394(196) ; 4396(225)
g73 not 4393(195) ; 4121(228)
g74 not 3749(194) ; 3751(229)
g75 not 3743(193) ; 3745(231)
g76 not 3737(192) ; 3739(233)
g77 not 3729(191) ; 3731(235)
g78 not 3723(190) ; 3725(237)
g79 not 3717(189) ; 3719(239)
g80 not 3711(188) ; 3713(241)
g81 not 3705(187) ; 3707(243)
g82 not 3701(186) ; 3703(245)
g83 not 3698(185) ; 3700(247)
g84 not 2256(184) ; 2258(249)
g85 not 2256(184) ; 1192(251)
g86 not 2253(183) ; 2255(252)
g87 not 2253(183) ; 1186(254)
g88 not 2247(182) ; 2249(255)
g89 not 2239(181) ; 2241(257)
g90 not 2236(180) ; 2238(259)
g91 not 2236(180) ; 1178(261)
g92 not 2230(179) ; 2232(262)
g93 not 2224(178) ; 2226(264)
g94 not 2218(177) ; 2220(266)
g95 not 2211(176) ; 2213(268)
g96 not 2208(175) ; 2210(270)
g97 not 2204(174) ; 2207(272)
g98 not 1496(173) ; 1499(273)
g99 or 1496(173)* 4528(206)* ; 1541(275)
g100 not 1492(172) ; 1495(276)
g101 and 1492(172) 4528(206) ; 1518(278)
g102 not 1486(171) ; 1488(279)
g103 not 1480(170) ; 1482(281)
g104 not 1469(169) ; 1471(283)
g105 not 1462(168) ; 1464(285)
g106 not 1459(167) ; 1461(287)
g107 not 1455(166) ; 1458(289)
g108 and 186(109) 185(108) 182(105) 183(106) ; 4442(290)
g109 and 199(122) 188(111) 172(95) 162(85) ; 1501(291)
g110 and 230(153) 218(141) 152(75) 210(133) ; 4514(292)
g111 and 240(163) 228(151) 184(107) 150(73) ; 2857(293)
g112 and 133(66) 134(67) ; 1184(294)
g113 and 106(53) ; 446(393)
g114 not 106(53) ; 1500(296)
g115 not 57(20) ; 400(297)
g116 and 38(11) ; 1210(298)
g117 and 38(11) ; 1198(299)
g118 and 18(5) ; 1512(300)
g119 and 18(5) ; 1524(301)
g120 not 18(5) ; 1535(302)
g121 and 18(5) ; 1503(303)
g122 and 15(4) ; 1205(305)
g123 or 9(2)* 12(3)* ; 1206(306)
g124 or 9(2)* 12(3)* ; 1207(307)
g125 not 5(1) ; 574(308)
g126 not 5(1) ; 575(309)
g127 not 5(1) ; 401(310)
g128 and 1(0) ; 432(428)
g129 or 2207(272)* 4528(206)* ; 2883(314)
g130 and 1458(289) 4528(206) ; 2871(315)
g131 not 4833(207) ; 4839(316)
g132 not 2828(208) ; 2833(317)
g133 and 4439(209) ; 6853(318)
g134 and 4439(209) ; 6567(319)
g135 and 4434(211) ; 6575(320)
g136 and 4434(211) ; 6861(321)
g137 and 4429(213) ; 6583(322)
g138 and 4429(213) ; 6869(323)
g139 and 4422(215) ; 6909(324)
g140 and 4422(215) ; 6591(325)
g141 and 4417(217) ; 6877(326)
g142 and 4417(217) ; 6599(327)
g143 and 4412(219) ; 6607(328)
g144 and 4412(219) ; 6885(329)
g145 and 4407(221) ; 6893(330)
g146 and 4407(221) ; 6615(331)
g147 and 4402(223) ; 6901(332)
g148 and 4402(223) ; 6623(333)
g149 and 4396(225) ; 6631(334)
g150 and 4396(225) ; 6917(335)
g151 and 3751(229) ; 5985(336)
g152 and 3751(229) ; 5865(337)
g153 and 3745(231) ; 5873(338)
g154 and 3745(231) ; 5993(339)
g155 and 3739(233) ; 6001(340)
g156 and 3739(233) ; 5881(341)
g157 and 3731(235) ; 6041(342)
g158 and 3731(235) ; 5889(343)
g159 and 3725(237) ; 5897(344)
g160 and 3725(237) ; 6009(345)
g161 and 3719(239) ; 6017(346)
g162 and 3719(239) ; 5905(347)
g163 and 3713(241) ; 5913(348)
g164 and 3713(241) ; 6025(349)
g165 and 3707(243) ; 6033(350)
g166 and 3707(243) ; 5921(351)
g167 and 1192(251) ; 5393(352)
g168 and 1192(251) ; 5745(353)
g169 and 1186(254) ; 5753(354)
g170 and 1186(254) ; 5401(355)
g171 and 2249(255) ; 5409(356)
g172 and 2249(255) ; 5761(357)
g173 and 2241(257) ; 5769(358)
g174 and 2241(257) ; 5449(359)
g175 and 1178(261) ; 5417(360)
g176 and 1178(261) ; 5777(361)
g177 and 2232(262) ; 5785(362)
g178 and 2232(262) ; 5425(363)
g179 and 2226(264) ; 5433(364)
g180 and 2226(264) ; 5793(365)
g181 and 2220(266) ; 5801(366)
g182 and 2220(266) ; 5441(367)
g183 and 2213(268) ; 5457(368)
g184 and 2213(268) ; 5809(369)
g185 and 1198(299) 1541(275) ; 777(370)
g186 and 1198(299) 1541(275) ; 1115(371)
g187 and 1541(275) ; 5175(372)
g188 and 1541(275) ; 4873(373)
g189 not 1518(278) ; 1519(374)
g190 and 1488(279) ; 4881(375)
g191 and 1488(279) ; 5191(376)
g192 and 1482(281) ; 5199(377)
g193 and 1482(281) ; 4889(378)
g194 and 1471(283) ; 5215(379)
g195 and 1471(283) ; 4905(380)
g196 and 1464(285) ; 4921(381)
g197 and 1464(285) ; 5223(382)
g198 and 1501(291) 4442(290) ; 2878(386)
g199 and 4514(292) 2857(293) ; 2876(389)
g200 and 575(309) 1184(294) ; 280(391)
g201 not 446(393) ; 1477(394)
g202 and 1210(298) ; 6554(396)
g203 and 1210(298) ; 6514(397)
g204 and 1198(299) ; 5186(398)
g205 and 1198(299) ; 5178(399)
g206 and 1198(299) ; 4916(400)
g207 and 1198(299) ; 4876(401)
g208 and 1512(300) ; 587(402)
g209 and 1512(300) ; 606(403)
g210 and 1512(300) ; 657(404)
g211 and 1512(300) ; 1336(405)
g212 not 1512(300) ; 1514(406)
g213 and 1524(301) ; 3622(407)
g214 and 1524(301) ; 3635(408)
g215 and 1524(301) ; 4640(409)
g216 and 1524(301) ; 4653(410)
g217 not 1524(301) ; 1530(411)
g218 and 1535(302) ; 3755(412)
g219 and 1535(302) ; 2259(413)
g220 and 1503(303) ; 678(414)
g221 and 1503(303) ; 1350(415)
g222 and 1503(303) ; 2892(416)
g223 and 1503(303) ; 2909(417)
g224 not 1503(303) ; 1507(418)
g225 and 1206(306) ; 581(421)
g226 and 1206(306) ; 601(422)
g227 and 1206(306) ; 650(423)
g228 and 1207(307) ; 671(424)
g229 and 1207(307) ; 2886(425)
g230 and 1207(307) ; 2905(426)
g231 and 432(428) ; 453(596)
g232 and 2883(314) ; 6511(429)
g233 not 2871(315) ; 2872(430)
g234 not 6853(318) ; 6859(431)
g235 not 6567(319) ; 6573(432)
g236 not 6575(320) ; 6581(433)
g237 not 6861(321) ; 6867(434)
g238 not 6583(322) ; 6589(435)
g239 not 6869(323) ; 6875(436)
g240 not 6909(324) ; 6915(437)
g241 not 6591(325) ; 6597(438)
g242 not 6877(326) ; 6883(439)
g243 not 6599(327) ; 6605(440)
g244 not 6607(328) ; 6613(441)
g245 not 6885(329) ; 6891(442)
g246 not 6893(330) ; 6899(443)
g247 not 6615(331) ; 6621(444)
g248 not 6901(332) ; 6907(445)
g249 not 6623(333) ; 6629(446)
g250 not 6631(334) ; 6637(447)
g251 not 6917(335) ; 6923(448)
g252 not 5985(336) ; 5991(449)
g253 not 5865(337) ; 5871(450)
g254 not 5873(338) ; 5879(451)
g255 not 5993(339) ; 5999(452)
g256 not 6001(340) ; 6007(453)
g257 not 5881(341) ; 5887(454)
g258 not 6041(342) ; 6047(455)
g259 not 5889(343) ; 5895(456)
g260 not 5897(344) ; 5903(457)
g261 not 6009(345) ; 6015(458)
g262 not 6017(346) ; 6023(459)
g263 not 5905(347) ; 5911(460)
g264 not 5913(348) ; 5919(461)
g265 not 6025(349) ; 6031(462)
g266 not 6033(350) ; 6039(463)
g267 not 5921(351) ; 5927(464)
g268 and 4653(410) 2258(249) ; 4685(465)
g269 not 5393(352) ; 5399(466)
g270 not 5745(353) ; 5751(467)
g271 and 4653(410) 2255(252) ; 4683(468)
g272 not 5753(354) ; 5759(469)
g273 not 5401(355) ; 5407(470)
g274 and 4653(410) 2249(255) ; 4681(471)
g275 not 5409(356) ; 5415(472)
g276 not 5761(357) ; 5767(473)
g277 not 5769(358) ; 5775(474)
g278 not 5449(359) ; 5455(475)
g279 and 4653(410) 2241(257) ; 4679(476)
g280 and 4653(410) 2238(259) ; 4677(477)
g281 not 5417(360) ; 5423(478)
g282 not 5777(361) ; 5783(479)
g283 not 5785(362) ; 5791(480)
g284 not 5425(363) ; 5431(481)
g285 and 4640(409) 2232(262) ; 4675(482)
g286 and 4640(409) 2226(264) ; 4673(483)
g287 not 5433(364) ; 5439(484)
g288 not 5793(365) ; 5799(485)
g289 not 5801(366) ; 5807(486)
g290 not 5441(367) ; 5447(487)
g291 and 4640(409) 2220(266) ; 4671(488)
g292 not 5457(368) ; 5463(489)
g293 and 4640(409) 2213(268) ; 4669(490)
g294 not 5809(369) ; 5815(491)
g295 and 4640(409) 2210(270) ; 4667(492)
g296 and 3635(408) 1499(273) ; 3663(493)
g297 not 5175(372) ; 5181(494)
g298 not 4873(373) ; 4879(495)
g299 and 3635(408) 1495(276) ; 3661(496)
g300 and 1519(374) ; 4913(497)
g301 and 1519(374) ; 5183(498)
g302 and 3635(408) 1488(279) ; 3659(499)
g303 not 4881(375) ; 4887(500)
g304 not 5191(376) ; 5197(501)
g305 not 5199(377) ; 5205(502)
g306 not 4889(378) ; 4895(503)
g307 and 3622(407) 1482(281) ; 3657(504)
g308 not 5215(379) ; 5221(505)
g309 and 3622(407) 1471(283) ; 3653(506)
g310 not 4905(380) ; 4911(507)
g311 not 4921(381) ; 4927(508)
g312 and 3622(407) 1464(285) ; 3651(509)
g313 not 5223(382) ; 5229(510)
g314 and 3622(407) 1461(287) ; 3649(511)
g315 and 2892(416) 216(139) ; 2921(512)
g316 and 2892(416) 215(138) ; 2923(513)
g317 and 2892(416) 214(137) ; 2925(514)
g318 and 2909(417) 213(136) ; 2927(515)
g319 and 2909(417) 212(135) ; 2929(516)
g320 and 2909(417) 211(134) ; 2931(517)
g321 and 2892(416) 209(132) ; 2919(518)
g322 and 1336(405) 181(104) ; 1364(519)
g323 and 1336(405) 180(103) ; 1368(520)
g324 and 1336(405) 179(102) ; 1370(521)
g325 and 1336(405) 178(101) ; 1372(522)
g326 and 657(404) 177(100) ; 691(523)
g327 and 657(404) 176(99) ; 693(524)
g328 and 657(404) 175(98) ; 695(525)
g329 and 657(404) 174(97) ; 697(526)
g330 and 657(404) 173(96) ; 699(527)
g331 and 1336(405) 171(94) ; 1366(528)
g332 and 587(402) 170(93) ; 615(529)
g333 and 587(402) 169(92) ; 617(530)
g334 and 587(402) 168(91) ; 619(531)
g335 and 587(402) 167(90) ; 621(532)
g336 and 606(403) 166(89) ; 623(533)
g337 and 606(403) 165(88) ; 625(534)
g338 and 606(403) 164(87) ; 627(535)
g339 and 1350(415) 161(84) ; 1374(537)
g340 and 1350(415) 160(83) ; 1378(538)
g341 and 1350(415) 159(82) ; 1380(539)
g342 and 1350(415) 158(81) ; 1382(540)
g343 and 678(414) 157(80) ; 701(541)
g344 and 678(414) 156(79) ; 703(542)
g345 and 678(414) 155(78) ; 705(543)
g346 and 678(414) 154(77) ; 707(544)
g347 and 678(414) 153(76) ; 709(545)
g348 and 1350(415) 151(74) ; 1376(546)
g349 and 1477(394) ; 4897(548)
g350 and 1477(394) ; 5207(549)
g351 and 3622(407) 1500(296) ; 3655(550)
g352 and 3755(412) 66(29) ; 3790(551)
g353 and 3755(412) 50(15) ; 3788(552)
g354 and 3755(412) 47(14) ; 3782(553)
g355 and 2259(413) 44(13) ; 2286(554)
g356 and 2259(413) 41(12) ; 2288(555)
g357 not 6554(396) ; 6558(556)
g358 and 1210(298) 2883(314) ; 3221(557)
g359 not 6514(397) ; 6518(558)
g360 and 1198(299) 1519(374) ; 784(559)
g361 and 1519(374) 1198(299) ; 1014(560)
g362 and 1519(374)* 1198(299)* ; 5231(561)
g363 not 5186(398) ; 5190(562)
g364 not 5178(399) ; 5182(563)
g365 and 1198(299)* 1519(374)* ; 4929(564)
g366 not 4916(400) ; 4920(565)
g367 not 4876(401) ; 4880(566)
g368 and 3755(412) 35(10) ; 3784(567)
g369 and 3755(412) 32(9) ; 3786(568)
g370 and 2259(413) 29(8) ; 2290(569)
g371 and 2259(413) 26(7) ; 2292(570)
g372 and 2259(413) 23(6) ; 2294(571)
g373 not 587(402) ; 594(572)
g374 not 606(403) ; 611(573)
g375 not 657(404) ; 664(574)
g376 not 1336(405) ; 1343(575)
g377 and 1514(406) ; 2019(576)
g378 and 1514(406) ; 2117(577)
g379 not 3622(407) ; 3629(578)
g380 not 3635(408) ; 3642(579)
g381 not 4640(409) ; 4647(580)
g382 not 4653(410) ; 4660(581)
g383 and 1530(411) ; 4444(582)
g384 and 1530(411) ; 4457(583)
g385 and 1530(411) ; 4094(584)
g386 and 1530(411) ; 4107(585)
g387 not 3755(412) ; 3762(586)
g388 not 2259(413) ; 2266(587)
g389 not 678(414) ; 685(588)
g390 not 1350(415) ; 1357(589)
g391 not 2892(416) ; 2899(590)
g392 not 2909(417) ; 2914(591)
g393 and 1507(418) ; 2032(592)
g394 and 1507(418) ; 2130(593)
g395 and 1507(418) ; 2272(594)
g396 and 1507(418) ; 3768(595)
g397 or 6518(558)* 6511(429)* ; 3169(597)
g398 not 6511(429) ; 6517(598)
g399 and 2872(430) ; 6551(599)
g400 and 3642(579) 3703(245) ; 3665(600)
g401 and 3642(579) 2204(174) ; 3662(601)
g402 or 5182(563)* 5175(372)* ; 1006(602)
g403 or 4880(566)* 4873(373)* ; 764(603)
g404 or 4920(565)* 4913(497)* ; 886(604)
g405 not 4913(497) ; 4919(605)
g406 or 5190(562)* 5183(498)* ; 1018(606)
g407 not 5183(498) ; 5189(607)
g408 and 3642(579) 1455(166) ; 3660(608)
g409 or 2921(512) 2899(590) ; 2922(609)
g410 or 2923(513) 2899(590) ; 2924(610)
g411 or 2925(514) 2899(590) ; 2926(611)
g412 or 2927(515) 2914(591) ; 2928(612)
g413 or 2929(516) 2914(591) ; 2930(613)
g414 or 2931(517) 2914(591) ; 2932(614)
g415 or 2919(518) 2899(590) ; 2920(615)
g416 and 2266(587) 208(131) ; 2285(616)
g417 and 2266(587) 207(130) ; 2289(617)
g418 and 2266(587) 206(129) ; 2291(618)
g419 and 2266(587) 205(128) ; 2293(619)
g420 and 2266(587) 198(121) ; 2287(620)
g421 and 3762(586) 193(116) ; 3781(621)
g422 and 3762(586) 192(115) ; 3783(622)
g423 and 3762(586) 191(114) ; 3785(623)
g424 and 3762(586) 190(113) ; 3787(624)
g425 and 3762(586) 189(112) ; 3789(625)
g426 or 691(523) 664(574) ; 692(626)
g427 or 693(524) 664(574) ; 694(627)
g428 or 695(525) 664(574) ; 696(628)
g429 or 697(526) 664(574) ; 698(629)
g430 or 699(527) 664(574) ; 700(630)
g431 or 615(529) 594(572) ; 577(631)
g432 or 617(530) 594(572) ; 618(632)
g433 or 619(531) 594(572) ; 620(633)
g434 or 621(532) 594(572) ; 622(634)
g435 or 623(533) 611(573) ; 624(635)
g436 or 625(534) 611(573) ; 626(636)
g437 or 627(535) 611(573) ; 628(637)
g438 or 701(541) 685(588) ; 702(638)
g439 or 703(542) 685(588) ; 704(639)
g440 or 705(543) 685(588) ; 706(640)
g441 or 707(544) 685(588) ; 708(641)
g442 or 709(545) 685(588) ; 710(642)
g443 and 1357(589) 147(72) ; 1375(643)
g444 and 1343(575) 147(72) ; 1365(644)
g445 and 1357(589) 144(71) ; 1379(645)
g446 and 1343(575) 144(71) ; 1369(646)
g447 and 1343(575) 141(70) ; 1363(647)
g448 and 1357(589) 141(70) ; 1373(648)
g449 and 1357(589) 138(69) ; 1377(649)
g450 and 1343(575) 138(69) ; 1367(650)
g451 and 1357(589) 135(68) ; 1381(651)
g452 and 1343(575) 135(68) ; 1371(652)
g453 and 2019(576) 130(65) ; 2048(653)
g454 and 2032(592) 130(65) ; 2058(654)
g455 and 2032(592) 127(64) ; 2060(655)
g456 and 2019(576) 127(64) ; 2050(656)
g457 and 2032(592) 124(63) ; 2062(657)
g458 and 2019(576) 124(63) ; 2052(658)
g459 and 2130(593) 121(62) ; 2162(659)
g460 and 2117(577) 121(62) ; 2152(660)
g461 and 2117(577) 118(61) ; 2146(661)
g462 and 2130(593) 118(61) ; 2156(662)
g463 and 2117(577) 115(60) ; 2144(663)
g464 and 2130(593) 115(60) ; 2154(664)
g465 and 3629(578) 114(59) ; 3648(665)
g466 and 3629(578) 113(58) ; 3650(666)
g467 and 3629(578) 112(57) ; 3656(667)
g468 and 3629(578) 111(56) ; 3652(668)
g469 and 4660(581) 110(55) ; 4684(669)
g470 and 4660(581) 109(54) ; 4682(670)
g471 not 4897(548) ; 4903(671)
g472 not 5207(549) ; 5213(672)
g473 and 2019(576) 103(52) ; 2046(673)
g474 and 2032(592) 103(52) ; 2056(674)
g475 and 2032(592) 100(51) ; 2064(675)
g476 and 2019(576) 100(51) ; 2054(676)
g477 and 2130(593) 97(50) ; 2158(677)
g478 and 2117(577) 97(50) ; 2148(678)
g479 and 2130(593) 94(49) ; 2160(679)
g480 and 2117(577) 94(49) ; 2150(680)
g481 and 3642(579) 88(47) ; 3658(681)
g482 and 3629(578) 87(46) ; 3654(682)
g483 and 4660(581) 86(45) ; 4680(683)
g484 and 4647(580) 85(44) ; 4674(684)
g485 and 4647(580) 84(43) ; 4672(685)
g486 and 4647(580) 83(42) ; 4670(686)
g487 and 4647(580) 82(41) ; 4666(687)
g488 and 4094(584) 81(40) ; 4135(688)
g489 and 4107(585) 80(39) ; 4138(689)
g490 and 4107(585) 79(38) ; 4141(690)
g491 and 4094(584) 78(37) ; 4129(691)
g492 and 4094(584) 77(36) ; 4126(692)
g493 and 4444(582) 76(35) ; 4477(693)
g494 and 4444(582) 75(34) ; 4479(694)
g495 and 4444(582) 74(33) ; 4475(695)
g496 and 4457(583) 73(32) ; 4481(696)
g497 and 4444(582) 70(31) ; 4473(697)
g498 and 3642(579) 70(31) ; 3666(698)
g499 and 4444(582) 69(30) ; 4471(699)
g500 and 3768(595) 66(29) ; 3800(700)
g501 and 4647(580) 65(28) ; 4668(701)
g502 and 4660(581) 64(27) ; 4676(702)
g503 and 4660(581) 63(26) ; 4678(703)
g504 and 4107(585) 62(25) ; 4150(704)
g505 and 4107(585) 61(24) ; 4147(705)
g506 and 4107(585) 60(23) ; 4144(706)
g507 and 4094(584) 59(22) ; 4132(707)
g508 and 4094(584) 58(21) ; 4123(708)
g509 and 4457(583) 56(19) ; 4489(709)
g510 and 4457(583) 55(18) ; 4487(710)
g511 and 4457(583) 54(17) ; 4485(711)
g512 and 4457(583) 53(16) ; 4483(712)
g513 and 3768(595) 50(15) ; 3798(713)
g514 and 3768(595) 47(14) ; 3792(714)
g515 and 2272(594) 44(13) ; 2296(715)
g516 and 2272(594) 41(12) ; 2298(716)
g517 and 1210(298) 2872(430) ; 3173(717)
g518 and 784(559) ; 4970(718)
g519 and 1014(560) ; 5239(719)
g520 not 5231(561) ; 5237(720)
g521 or 5181(494)* 5178(399)* ; 1005(721)
g522 not 4929(564) ; 4935(722)
g523 or 4879(495)* 4876(401)* ; 763(723)
g524 and 3768(595) 35(10) ; 3794(724)
g525 and 3768(595) 32(9) ; 3796(725)
g526 and 2272(594) 29(8) ; 2300(726)
g527 and 2272(594) 26(7) ; 2302(727)
g528 and 2272(594) 23(6) ; 2304(728)
g529 or 587(402) 594(572) ; 616(729)
g530 not 2019(576) ; 2026(730)
g531 not 2117(577) ; 2124(731)
g532 not 4444(582) ; 4451(732)
g533 not 4457(583) ; 4464(733)
g534 not 4094(584) ; 4101(734)
g535 not 4107(585) ; 4114(735)
g536 or 2892(416) 2899(590) ; 2918(736)
g537 not 2032(592) ; 2039(737)
g538 not 2130(593) ; 2137(738)
g539 not 2272(594) ; 2279(739)
g540 not 3768(595) ; 3775(740)
g541 not 6551(599) ; 6557(741)
g542 and 4114(735) 4439(209) ; 4149(742)
g543 and 4114(735) 4434(211) ; 4146(743)
g544 and 4114(735) 4429(213) ; 4143(744)
g545 and 4114(735) 4422(215) ; 4140(745)
g546 and 4114(735) 4417(217) ; 4137(746)
g547 and 4101(734) 4412(219) ; 4134(747)
g548 and 4101(734) 4407(221) ; 4131(748)
g549 and 4101(734) 4402(223) ; 4128(749)
g550 and 4101(734) 4396(225) ; 4125(750)
g551 and 4101(734) 4121(228) ; 4122(751)
g552 and 4464(733) 3751(229) ; 4488(752)
g553 and 4464(733) 3745(231) ; 4486(753)
g554 and 4464(733) 3739(233) ; 4484(754)
g555 and 4464(733) 3731(235) ; 4482(755)
g556 and 4464(733) 3725(237) ; 4480(756)
g557 and 4451(732) 3719(239) ; 4478(757)
g558 and 4451(732) 3713(241) ; 4476(758)
g559 and 4451(732) 3707(243) ; 4474(759)
g560 and 4451(732) 3703(245) ; 4472(760)
g561 and 4451(732) 3700(247) ; 4470(761)
g562 or 4685(465) 4684(669) ; 4710(762)
g563 or 4683(468) 4682(670) ; 4707(763)
g564 or 4681(471) 4680(683) ; 4704(764)
g565 or 4679(476) 4678(703) ; 4701(765)
g566 or 4677(477) 4676(702) ; 4698(766)
g567 or 4675(482) 4674(684) ; 4695(767)
g568 or 4673(483) 4672(685) ; 4692(768)
g569 or 4671(488) 4670(686) ; 4689(769)
g570 or 4669(490) 4668(701) ; 4686(770)
g571 or 4667(492) 4666(687) ; 7466(771)
g572 or 3663(493) 3662(601) ; 6711(772)
g573 or 1006(602)* 1005(721)* ; 1007(773)
g574 or 764(603)* 763(723)* ; 765(774)
g575 or 3661(496) 3660(608) ; 6714(775)
g576 or 3659(499) 3658(681) ; 3679(776)
g577 or 3657(504) 3656(667) ; 3676(777)
g578 or 3653(506) 3652(668) ; 3670(778)
g579 or 3651(509) 3650(666) ; 3667(779)
g580 or 3649(511) 3648(665) ; 6690(780)
g581 and 2279(739) 239(162) ; 2295(781)
g582 and 2279(739) 238(161) ; 2299(782)
g583 and 2279(739) 237(160) ; 2301(783)
g584 and 2279(739) 236(159) ; 2303(784)
g585 and 2039(737) 235(158) ; 2055(785)
g586 and 2039(737) 234(157) ; 2057(786)
g587 and 2039(737) 233(156) ; 2059(787)
g588 and 2039(737) 232(155) ; 2061(788)
g589 and 2039(737) 231(154) ; 2063(789)
g590 and 2279(739) 229(152) ; 2297(790)
g591 and 2137(738) 227(150) ; 2153(791)
g592 and 2137(738) 226(149) ; 2157(792)
g593 and 2137(738) 225(148) ; 2159(793)
g594 and 2137(738) 224(147) ; 2161(794)
g595 and 3775(740) 223(146) ; 3791(795)
g596 and 3775(740) 222(145) ; 3793(796)
g597 and 3775(740) 221(144) ; 3795(797)
g598 and 3775(740) 220(143) ; 3797(798)
g599 and 3775(740) 219(142) ; 3799(799)
g600 and 2137(738) 217(140) ; 2155(800)
g601 and 2026(730) 204(127) ; 2045(801)
g602 and 2026(730) 203(126) ; 2047(802)
g603 and 2026(730) 202(125) ; 2049(803)
g604 and 2026(730) 201(124) ; 2051(804)
g605 and 2026(730) 200(123) ; 2053(805)
g606 and 2124(731) 197(120) ; 2143(806)
g607 and 2124(731) 196(119) ; 2147(807)
g608 and 2124(731) 195(118) ; 2149(808)
g609 and 2124(731) 194(117) ; 2151(809)
g610 and 2124(731) 187(110) ; 2145(810)
g611 or 1364(519) 1363(647) ; 7296(811)
g612 or 1368(520) 1367(650) ; 1387(812)
g613 or 1370(521) 1369(646) ; 1391(813)
g614 or 1372(522) 1371(652) ; 1395(814)
g615 or 1366(528) 1365(644) ; 1383(815)
g616 or 1374(537) 1373(648) ; 5318(816)
g617 or 1378(538) 1377(649) ; 1406(817)
g618 or 1380(539) 1379(645) ; 1412(818)
g619 or 1382(540) 1381(651) ; 1418(819)
g620 or 1376(546) 1375(643) ; 1399(820)
g621 or 3655(550) 3654(682) ; 3673(821)
g622 or 3790(551) 3789(625) ; 3813(822)
g623 or 3788(552) 3787(624) ; 3810(823)
g624 or 3782(553) 3781(621) ; 3801(824)
g625 or 2286(554) 2285(616) ; 7252(825)
g626 or 2288(555) 2287(620) ; 2305(826)
g627 or 6558(556)* 6551(599)* ; 3211(827)
g628 or 6517(598)* 6514(397)* ; 3168(828)
g629 not 4970(718) ; 4976(829)
g630 not 5239(719) ; 5245(830)
g631 or 5189(607)* 5186(398)* ; 1017(831)
g632 or 4919(605)* 4916(400)* ; 885(832)
g633 or 3784(567) 3783(622) ; 3804(833)
g634 or 3786(568) 3785(623) ; 3807(834)
g635 or 2290(569) 2289(617) ; 2308(835)
g636 or 2292(570) 2291(618) ; 2312(836)
g637 or 2294(571) 2293(619) ; 2316(837)
g638 or 3635(408) 3666(698) ; 3686(838)
g639 or 3635(408) 3665(600) ; 3682(839)
g640 and 581(421) 577(631) ; 579(840)
g641 and 581(421) 622(634) ; 641(841)
g642 and 581(421) 620(633) ; 637(842)
g643 and 581(421) 618(632) ; 633(843)
g644 and 581(421) 616(729) ; 629(844)
g645 and 601(422) 628(637) ; 5305(845)
g646 and 601(422) 626(636) ; 5308(846)
g647 and 601(422) 624(635) ; 645(847)
g648 and 650(423) 700(630) ; 727(848)
g649 and 650(423) 698(629) ; 723(849)
g650 and 650(423) 696(628) ; 719(850)
g651 and 650(423) 694(627) ; 715(851)
g652 and 650(423) 692(626) ; 711(852)
g653 and 671(424) 706(640) ; 745(853)
g654 and 671(424) 704(639) ; 737(854)
g655 and 671(424) 702(638) ; 731(855)
g656 and 671(424) 710(642) ; 757(856)
g657 and 671(424) 708(641) ; 751(857)
g658 and 2886(425) 2926(611) ; 2946(858)
g659 and 2886(425) 2924(610) ; 2942(859)
g660 and 2886(425) 2922(609) ; 2938(860)
g661 and 2886(425) 2920(615) ; 2933(861)
g662 and 2886(425) 2918(736) ; 4525(862)
g663 and 2905(426) 2932(614) ; 5271(863)
g664 and 2905(426) 2930(613) ; 5274(864)
g665 and 2905(426) 2928(612) ; 2950(865)
g666 or 3169(597)* 3168(828)* ; 3170(866)
g667 and 727(848) 4710(762) ; 2962(867)
g668 and 4710(762) ; 7497(868)
g669 and 4710(762) ; 6367(869)
g670 and 757(856) 1192(251) ; 1553(870)
g671 and 757(856) 1192(251) ; 1802(871)
g672 and 723(849) 4707(763) ; 2970(872)
g673 and 4707(763) ; 7500(873)
g674 and 4707(763) ; 6375(874)
g675 and 751(857) 1186(254) ; 1816(875)
g676 and 751(857) 1186(254) ; 1567(876)
g677 and 745(853) 2249(255) ; 1584(877)
g678 and 745(853) 2249(255) ; 1834(878)
g679 and 719(850) 4704(764) ; 2977(879)
g680 and 4704(764) ; 6383(880)
g681 and 4704(764) ; 7487(881)
g682 and 737(854) 2241(257) ; 1590(882)
g683 and 2241(257) 737(854) ; 1841(883)
g684 and 2241(257)* 737(854)* ; 5849(884)
g685 and 737(854)* 2241(257)* ; 5465(885)
g686 and 715(851) 4701(765) ; 2979(886)
g687 and 4701(765) ; 7490(887)
g688 and 4701(765) ; 6423(888)
g689 and 711(852) 4698(766) ; 2989(889)
g690 and 4698(766) ; 7479(890)
g691 and 4698(766) ; 6391(891)
g692 and 731(855) 1178(261) ; 1606(892)
g693 and 731(855) 1178(261) ; 1866(893)
g694 and 1418(819) 2232(262) ; 1624(894)
g695 and 1418(819) 2232(262) ; 1880(895)
g696 and 1395(814) 4695(767) ; 2998(896)
g697 and 4695(767) ; 6399(897)
g698 and 4695(767) ; 7482(898)
g699 and 1412(818) 2226(264) ; 1647(899)
g700 and 1412(818) 2226(264) ; 1897(900)
g701 and 1391(813) 4692(768) ; 3006(901)
g702 and 4692(768) ; 7471(902)
g703 and 4692(768) ; 6407(903)
g704 and 1406(817) 2220(266) ; 1669(904)
g705 and 1406(817) 2220(266) ; 1914(905)
g706 and 1387(812) 4689(769) ; 3013(906)
g707 and 4689(769) ; 6415(907)
g708 and 4689(769) ; 7474(908)
g709 and 1399(820) 2213(268) ; 1677(909)
g710 and 1399(820) 2213(268) ; 1929(910)
g711 and 1399(820)* 2213(268)* ; 5581(911)
g712 and 1383(815) 4686(770) ; 3015(912)
g713 and 4686(770) ; 7463(913)
g714 and 4686(770) ; 6431(914)
g715 not 7466(771) ; 7470(915)
g716 not 6711(772) ; 6717(916)
g717 and 1007(773) ; 5242(917)
g718 and 1007(773) ; 5234(918)
g719 and 765(774) ; 4962(919)
g720 and 765(774) ; 5003(920)
g721 not 6714(775) ; 6718(921)
g722 or 886(604)* 885(832)* ; 887(922)
g723 or 1018(606)* 1017(831)* ; 1019(923)
g724 and 2950(865) 1488(279) ; 802(924)
g725 and 2950(865) 1488(279) ; 1035(925)
g726 and 645(847) 3679(776) ; 3183(926)
g727 and 3679(776) ; 6703(927)
g728 and 3679(776) ; 6519(928)
g729 and 2946(858) 1482(281) ; 821(929)
g730 and 2946(858) 1482(281) ; 1050(930)
g731 and 641(841) 3676(777) ; 3192(931)
g732 and 3676(777) ; 6527(932)
g733 and 3676(777) ; 6706(933)
g734 and 2938(860) 1471(283) ; 868(934)
g735 and 2938(860) 1471(283) ; 1086(935)
g736 and 633(843) 3670(778) ; 3207(936)
g737 and 3670(778) ; 6543(937)
g738 and 3670(778) ; 6698(938)
g739 and 2933(861) 1464(285) ; 877(939)
g740 and 2933(861) 1464(285) ; 1102(940)
g741 and 2933(861)* 1464(285)* ; 5011(941)
g742 and 629(844) 3667(779) ; 3209(942)
g743 and 3667(779) ; 6687(943)
g744 and 3667(779) ; 6559(944)
g745 not 6690(780) ; 6694(945)
g746 not 7296(811) ; 7300(946)
g747 and 1387(812) ; 6418(947)
g748 and 1387(812) ; 7304(948)
g749 and 1391(813) ; 7301(949)
g750 and 1391(813) ; 6410(950)
g751 and 1395(814) ; 6402(951)
g752 and 1395(814) ; 7312(952)
g753 and 1383(815) ; 7293(953)
g754 and 1383(815) ; 6434(954)
g755 not 5318(816) ; 5322(955)
g756 and 1406(817) ; 5326(956)
g757 and 1406(817) ; 5444(957)
g758 and 1406(817) ; 5804(958)
g759 and 1412(818) ; 5323(959)
g760 and 1412(818) ; 5796(960)
g761 and 1412(818) ; 5436(961)
g762 and 1418(819) ; 5334(962)
g763 and 1418(819) ; 5428(963)
g764 and 1418(819) ; 5788(964)
g765 and 1399(820) ; 5315(965)
g766 and 1399(820) ; 5812(966)
g767 and 1399(820) ; 5460(967)
g768 or 2048(653) 2047(802) ; 2069(968)
g769 or 2058(654) 2057(786) ; 2091(969)
g770 or 2060(655) 2059(787) ; 2099(970)
g771 or 2050(656) 2049(803) ; 2073(971)
g772 or 2062(657) 2061(788) ; 2105(972)
g773 or 2052(658) 2051(804) ; 2077(973)
g774 or 2162(659) 2161(794) ; 2198(974)
g775 or 2152(660) 2151(809) ; 2175(975)
g776 or 2146(661) 2145(810) ; 2163(976)
g777 or 2156(662) 2155(800) ; 2179(977)
g778 or 2144(663) 2143(806) ; 7208(978)
g779 or 2154(664) 2153(791) ; 6724(979)
g780 and 2942(859) 1477(394) ; 845(980)
g781 and 2942(859) 1477(394) ; 1068(981)
g782 and 637(842) 3673(821) ; 3200(982)
g783 and 3673(821) ; 6695(983)
g784 and 3673(821) ; 6535(984)
g785 or 2046(673) 2045(801) ; 2065(985)
g786 or 2056(674) 2055(785) ; 2085(986)
g787 or 2064(675) 2063(789) ; 2111(987)
g788 or 2054(676) 2053(805) ; 2081(988)
g789 or 2158(677) 2157(792) ; 2186(989)
g790 or 2148(678) 2147(807) ; 2167(990)
g791 or 2160(679) 2159(793) ; 2192(991)
g792 or 2150(680) 2149(808) ; 2171(992)
g793 or 4135(688) 4134(747) ; 4160(993)
g794 or 4138(689) 4137(746) ; 4163(994)
g795 or 4141(690) 4140(745) ; 4166(995)
g796 or 4129(691) 4128(749) ; 4154(996)
g797 or 4126(692) 4125(750) ; 4151(997)
g798 or 4477(693) 4476(758) ; 4493(998)
g799 or 4479(694) 4478(757) ; 4496(999)
g800 or 4475(695) 4474(759) ; 4490(1000)
g801 or 4481(696) 4480(756) ; 4499(1001)
g802 or 4473(697) 4472(760) ; 7507(1002)
g803 or 4471(699) 4470(761) ; 7510(1003)
g804 or 3800(700) 3799(799) ; 3838(1004)
g805 and 3813(822) ; 7239(1005)
g806 and 3813(822) ; 6442(1006)
g807 or 4150(704) 4149(742) ; 4175(1007)
g808 or 4147(705) 4146(743) ; 4172(1008)
g809 or 4144(706) 4143(744) ; 4169(1009)
g810 or 4132(707) 4131(748) ; 4157(1010)
g811 or 4123(708) 4122(751) ; 7554(1011)
g812 or 4489(709) 4488(752) ; 4511(1012)
g813 or 4487(710) 4486(753) ; 4508(1013)
g814 or 4485(711) 4484(754) ; 4505(1014)
g815 or 4483(712) 4482(755) ; 4502(1015)
g816 or 3798(713) 3797(798) ; 3833(1016)
g817 and 3810(823) ; 6450(1017)
g818 and 3810(823) ; 7242(1018)
g819 and 3801(824) ; 6466(1019)
g820 and 3801(824) ; 7221(1020)
g821 or 3792(714) 3791(795) ; 3816(1021)
g822 not 7252(825) ; 7256(1022)
g823 or 2296(715) 2295(781) ; 6768(1023)
g824 and 2305(826) ; 7249(1024)
g825 or 2298(716) 2297(790) ; 2320(1025)
g826 or 6557(741)* 6554(396)* ; 3210(1026)
g827 and 784(559) 765(774) ; 913(1027)
g828 and 784(559) 765(774) ; 907(1028)
g829 and 784(559) 765(774) ; 915(1029)
g830 and 784(559) 765(774) ; 916(1030)
g831 and 1014(560) 1007(773) ; 1116(1031)
g832 and 3804(833) ; 6498(1032)
g833 and 3804(833) ; 7232(1033)
g834 or 3794(724) 3793(796) ; 3821(1034)
g835 or 3796(725) 3795(797) ; 3828(1035)
g836 and 3807(834) ; 6458(1036)
g837 and 3807(834) ; 7229(1037)
g838 or 2300(726) 2299(782) ; 2323(1038)
g839 and 2308(835) ; 7412(1039)
g840 and 2308(835) ; 7260(1040)
g841 or 2302(727) 2301(783) ; 2329(1041)
g842 and 2312(836) ; 7404(1042)
g843 and 2312(836) ; 7257(1043)
g844 or 2304(728) 2303(784) ; 2335(1044)
g845 and 2316(837) ; 7396(1045)
g846 and 2316(837) ; 7268(1046)
g847 and 3686(838) ; 7425(1047)
g848 and 3682(839) ; 5929(1048)
g849 and 3682(839) ; 6049(1049)
g850 and 2305(826) 1535(302) ; 3695(1050)
g851 not 579(840) ; 5284(1051)
g852 and 641(841) ; 5300(1052)
g853 and 641(841) ; 6530(1053)
g854 and 637(842) ; 5289(1054)
g855 and 637(842) ; 6538(1055)
g856 and 633(843) ; 5292(1056)
g857 and 633(843) ; 6546(1057)
g858 and 629(844) ; 5281(1058)
g859 and 629(844) ; 6562(1059)
g860 not 5305(845) ; 5311(1060)
g861 not 5308(846) ; 5312(1061)
g862 and 645(847) ; 5297(1062)
g863 and 645(847) ; 6522(1063)
g864 and 727(848) ; 7327(1064)
g865 and 727(848) ; 6370(1065)
g866 and 723(849) ; 6378(1066)
g867 and 723(849) ; 7330(1067)
g868 and 719(850) ; 7317(1068)
g869 and 719(850) ; 6386(1069)
g870 and 715(851) ; 6426(1070)
g871 and 715(851) ; 7320(1071)
g872 and 711(852) ; 7309(1072)
g873 and 711(852) ; 6394(1073)
g874 and 745(853) ; 5339(1074)
g875 and 745(853) ; 5764(1075)
g876 and 745(853) ; 5412(1076)
g877 and 737(854) ; 5452(1077)
g878 and 737(854) ; 5772(1078)
g879 and 737(854) ; 5342(1079)
g880 and 731(855) ; 5331(1080)
g881 and 731(855) ; 5780(1081)
g882 and 731(855) ; 5420(1082)
g883 and 757(856) ; 5349(1083)
g884 and 757(856) ; 5396(1084)
g885 and 757(856) ; 5748(1085)
g886 and 751(857) ; 5756(1086)
g887 and 751(857) ; 5404(1087)
g888 and 751(857) ; 5352(1088)
g889 and 2946(858) ; 5202(1089)
g890 and 2946(858) ; 4892(1090)
g891 and 2946(858) ; 5266(1091)
g892 and 2942(859) ; 5255(1092)
g893 and 2942(859) ; 4900(1093)
g894 and 2942(859) ; 5210(1094)
g895 and 2938(860) ; 5218(1095)
g896 and 2938(860) ; 4908(1096)
g897 and 2938(860) ; 5258(1097)
g898 and 2933(861) ; 5247(1098)
g899 and 2933(861) ; 4924(1099)
g900 and 2933(861) ; 5226(1100)
g901 not 4525(862) ; 5250(1101)
g902 not 5271(863) ; 5277(1102)
g903 not 5274(864) ; 5278(1103)
g904 and 2950(865) ; 5263(1104)
g905 and 2950(865) ; 4884(1105)
g906 and 2950(865) ; 5194(1106)
g907 and 3838(1004) 4439(209) ; 3292(1107)
g908 and 3838(1004) 4439(209) ; 3853(1108)
g909 and 3833(1016) 4434(211) ; 3308(1109)
g910 and 3833(1016) 4434(211) ; 3868(1110)
g911 and 3828(1035) 4429(213) ; 3327(1111)
g912 and 3828(1035) 4429(213) ; 3885(1112)
g913 and 4422(215) 3821(1034) ; 3335(1113)
g914 and 3821(1034) 4422(215) ; 3891(1114)
g915 and 3821(1034)* 4422(215)* ; 6925(1115)
g916 and 4422(215)* 3821(1034)* ; 6671(1116)
g917 and 3816(1021) 4417(217) ; 3362(1117)
g918 and 3816(1021) 4417(217) ; 3908(1118)
g919 and 2198(974) 4412(219) ; 3376(1119)
g920 and 2198(974) 4412(219) ; 3926(1120)
g921 and 2192(991) 4407(221) ; 3393(1121)
g922 and 2192(991) 4407(221) ; 3949(1122)
g923 and 2186(989) 4402(223) ; 3410(1123)
g924 and 2186(989) 4402(223) ; 3971(1124)
g925 and 2179(977) 4396(225) ; 3425(1125)
g926 and 2179(977) 4396(225) ; 3979(1126)
g927 and 2179(977)* 4396(225)* ; 7041(1127)
g928 and 2111(987) 3751(229) ; 2351(1128)
g929 and 2111(987) 3751(229) ; 2597(1129)
g930 and 2105(972) 3745(231) ; 2366(1130)
g931 and 2105(972) 3745(231) ; 2612(1131)
g932 and 2099(970) 3739(233) ; 2384(1132)
g933 and 2099(970) 3739(233) ; 2629(1133)
g934 and 3731(235) 2091(969) ; 2391(1134)
g935 and 2091(969) 3731(235) ; 2635(1135)
g936 and 2091(969)* 3731(235)* ; 6057(1136)
g937 and 3731(235)* 2091(969)* ; 5969(1137)
g938 and 2085(986) 3725(237) ; 2417(1138)
g939 and 2085(986) 3725(237) ; 2652(1139)
g940 and 2335(1044) 3719(239) ; 2431(1140)
g941 and 2335(1044) 3719(239) ; 2670(1141)
g942 and 2329(1041) 3713(241) ; 2448(1142)
g943 and 2329(1041) 3713(241) ; 2693(1143)
g944 and 2323(1038) 3707(243) ; 2465(1144)
g945 and 2323(1038) 3707(243) ; 2715(1145)
g946 not 7497(868) ; 7503(1146)
g947 not 6367(869) ; 6373(1147)
g948 or 5399(466)* 5396(1084)* ; 1544(1148)
g949 or 5751(467)* 5748(1085)* ; 1793(1149)
g950 not 7500(873) ; 7504(1150)
g951 not 6375(874) ; 6381(1151)
g952 or 5759(469)* 5756(1086)* ; 1803(1152)
g953 or 5407(470)* 5404(1087)* ; 1554(1153)
g954 not 6383(880) ; 6389(1154)
g955 not 7487(881) ; 7493(1155)
g956 or 5415(472)* 5412(1076)* ; 1571(1156)
g957 or 5767(473)* 5764(1075)* ; 1820(1157)
g958 and 1590(882) ; 5523(1158)
g959 and 1841(883) ; 5857(1159)
g960 or 5775(474)* 5772(1078)* ; 1848(1160)
g961 not 5849(884) ; 5855(1161)
g962 not 5465(885) ; 5471(1162)
g963 or 5455(475)* 5452(1077)* ; 1685(1163)
g964 not 7490(887) ; 7494(1164)
g965 not 6423(888) ; 6429(1165)
g966 not 7479(890) ; 7485(1166)
g967 not 6391(891) ; 6397(1167)
g968 or 5423(478)* 5420(1082)* ; 1596(1168)
g969 or 5783(479)* 5780(1081)* ; 1857(1169)
g970 or 5791(480)* 5788(964)* ; 1867(1170)
g971 or 5431(481)* 5428(963)* ; 1607(1171)
g972 not 6399(897) ; 6405(1172)
g973 not 7482(898) ; 7486(1173)
g974 not 7471(902) ; 7477(1174)
g975 not 6407(903) ; 6413(1175)
g976 or 5439(484)* 5436(961)* ; 1628(1176)
g977 or 5799(485)* 5796(960)* ; 1883(1177)
g978 or 5807(486)* 5804(958)* ; 1901(1178)
g979 or 5447(487)* 5444(957)* ; 1653(1179)
g980 not 6415(907) ; 6421(1180)
g981 not 7474(908) ; 7478(1181)
g982 and 1677(909) ; 5669(1182)
g983 not 5581(911) ; 5587(1183)
g984 or 5463(489)* 5460(967)* ; 1693(1184)
g985 or 7470(915)* 7463(913)* ; 4530(1185)
g986 not 7463(913) ; 7469(1186)
g987 not 6431(914) ; 6437(1187)
g988 or 5815(491)* 5812(966)* ; 1919(1188)
g989 or 6718(921)* 6711(772)* ; 6720(1189)
g990 or 916(1030) 777(370) ; 917(1190)
g991 and 915(1029)* 777(370)* ; 4983(1191)
g992 or 907(1028) 777(370) ; 908(1192)
g993 or 1116(1031) 1115(371) ; 1117(1193)
g994 not 5242(917) ; 5246(1194)
g995 not 5234(918) ; 5238(1195)
g996 and 1007(773) 1019(923) ; 1108(1196)
g997 and 765(774) 887(922) ; 953(1197)
g998 not 4962(919) ; 4966(1198)
g999 and 765(774) 887(922) ; 902(1199)
g1000 and 765(774) 887(922) ; 914(1200)
g1001 not 5003(920) ; 5007(1201)
g1002 or 6717(916)* 6714(775)* ; 6719(1202)
g1003 and 887(922) ; 4993(1203)
g1004 and 887(922) ; 4952(1204)
g1005 not 1019(923) ; 1023(1205)
g1006 not 6703(927) ; 6709(1206)
g1007 not 6519(928) ; 6525(1207)
g1008 or 4887(500)* 4884(1105)* ; 790(1208)
g1009 or 5197(501)* 5194(1106)* ; 1024(1209)
g1010 or 5205(502)* 5202(1089)* ; 1036(1210)
g1011 or 4895(503)* 4892(1090)* ; 803(1211)
g1012 not 6527(932) ; 6533(1212)
g1013 not 6706(933) ; 6710(1213)
g1014 or 5221(505)* 5218(1095)* ; 1072(1214)
g1015 not 6543(937) ; 6549(1215)
g1016 not 6698(938) ; 6702(1216)
g1017 or 4911(507)* 4908(1096)* ; 851(1217)
g1018 and 877(939) ; 5099(1218)
g1019 not 5011(941) ; 5017(1219)
g1020 or 4927(508)* 4924(1099)* ; 893(1220)
g1021 or 6694(945)* 6687(943)* ; 3503(1221)
g1022 not 6687(943) ; 6693(1222)
g1023 not 6559(944) ; 6565(1223)
g1024 or 5229(510)* 5226(1100)* ; 1091(1224)
g1025 or 7300(946)* 7293(953)* ; 4225(1225)
g1026 not 6418(947) ; 6422(1226)
g1027 not 7304(948) ; 7308(1227)
g1028 not 7301(949) ; 7307(1228)
g1029 not 6410(950) ; 6414(1229)
g1030 not 6402(951) ; 6406(1230)
g1031 not 7312(952) ; 7316(1231)
g1032 not 7293(953) ; 7299(1232)
g1033 not 6434(954) ; 6438(1233)
g1034 or 5322(955)* 5315(965)* ; 1262(1234)
g1035 not 5326(956) ; 5330(1235)
g1036 not 5444(957) ; 5448(1236)
g1037 not 5804(958) ; 5808(1237)
g1038 not 5323(959) ; 5329(1238)
g1039 not 5796(960) ; 5800(1239)
g1040 not 5436(961) ; 5440(1240)
g1041 not 5334(962) ; 5338(1241)
g1042 not 5428(963) ; 5432(1242)
g1043 not 5788(964) ; 5792(1243)
g1044 not 5315(965) ; 5321(1244)
g1045 not 5812(966) ; 5816(1245)
g1046 not 5460(967) ; 5464(1246)
g1047 and 2069(968) ; 7276(1247)
g1048 and 2069(968) 4502(1015) ; 4314(1248)
g1049 and 2069(968) ; 7420(1249)
g1050 and 2091(969) ; 5892(1250)
g1051 and 2091(969) ; 6044(1251)
g1052 and 2091(969) ; 6792(1252)
g1053 and 2099(970) ; 6789(1253)
g1054 and 2099(970) ; 6004(1254)
g1055 and 2099(970) ; 5884(1255)
g1056 and 2073(971) 4505(1014) ; 4312(1256)
g1057 and 2073(971) ; 7380(1257)
g1058 and 2073(971) ; 7273(1258)
g1059 and 2105(972) ; 5876(1259)
g1060 and 2105(972) ; 5996(1260)
g1061 and 2105(972) ; 6802(1261)
g1062 and 2077(973) 4508(1013) ; 4305(1262)
g1063 and 2077(973) ; 7372(1263)
g1064 and 2077(973) ; 7286(1264)
g1065 and 2198(974) ; 6740(1265)
g1066 and 2198(974) ; 6610(1266)
g1067 and 2198(974) ; 6888(1267)
g1068 and 2175(975) 4160(993) ; 3099(1268)
g1069 and 2175(975) ; 6474(1269)
g1070 and 2175(975) ; 7224(1270)
g1071 and 2163(976) 4151(997) ; 3116(1271)
g1072 and 2163(976) ; 6506(1272)
g1073 and 2163(976) ; 7205(1273)
g1074 and 2179(977) ; 6721(1274)
g1075 and 2179(977) ; 6634(1275)
g1076 and 2179(977) ; 6920(1276)
g1077 not 7208(978) ; 7212(1277)
g1078 not 6724(979) ; 6728(1278)
g1079 or 4903(671)* 4900(1093)* ; 825(1279)
g1080 or 5213(672)* 5210(1094)* ; 1053(1280)
g1081 not 6695(983) ; 6701(1281)
g1082 not 6535(984) ; 6541(1282)
g1083 and 2065(985) ; 7388(1283)
g1084 and 2065(985) 4499(1001) ; 4324(1284)
g1085 and 2065(985) ; 7265(1285)
g1086 and 2085(986) ; 6781(1286)
g1087 and 2085(986) ; 6012(1287)
g1088 and 2085(986) ; 5900(1288)
g1089 and 2111(987) ; 6799(1289)
g1090 and 2111(987) ; 5988(1290)
g1091 and 2111(987) ; 5868(1291)
g1092 and 2081(988) ; 7364(1292)
g1093 and 2081(988) 4511(1012) ; 4297(1293)
g1094 and 2081(988) ; 7283(1294)
g1095 and 2186(989) ; 6732(1295)
g1096 and 2186(989) ; 6904(1296)
g1097 and 2186(989) ; 6626(1297)
g1098 and 2167(990) 4154(996) ; 3114(1298)
g1099 and 2167(990) ; 6490(1299)
g1100 and 2167(990) ; 7216(1300)
g1101 and 2192(991) ; 6729(1301)
g1102 and 2192(991) ; 6896(1302)
g1103 and 2192(991) ; 6618(1303)
g1104 and 2171(992) ; 6482(1304)
g1105 and 2171(992) 4157(1010) ; 3107(1305)
g1106 and 2171(992) ; 7213(1306)
g1107 and 4160(993) ; 6471(1307)
g1108 and 4160(993) ; 7570(1308)
g1109 and 4163(994) ; 6463(1309)
g1110 and 4163(994) ; 7567(1310)
g1111 and 4166(995) ; 6495(1311)
g1112 and 4166(995) ; 7578(1312)
g1113 and 4154(996) ; 6487(1313)
g1114 and 4154(996) ; 7562(1314)
g1115 and 4151(997) ; 6503(1315)
g1116 and 4151(997) ; 7551(1316)
g1117 and 4493(998) ; 7515(1317)
g1118 and 4493(998) ; 7401(1318)
g1119 and 4496(999) ; 7393(1319)
g1120 and 4496(999) ; 7526(1320)
g1121 and 4490(1000) ; 7409(1321)
g1122 and 4490(1000) ; 7518(1322)
g1123 and 4499(1001) ; 7523(1323)
g1124 and 4499(1001) ; 7385(1324)
g1125 not 7507(1002) ; 7513(1325)
g1126 not 7510(1003) ; 7514(1326)
g1127 and 3838(1004) ; 6856(1327)
g1128 and 3838(1004) ; 6755(1328)
g1129 and 3838(1004) ; 6570(1329)
g1130 and 3813(822) 4175(1007) ; 3059(1330)
g1131 not 7239(1005) ; 7245(1331)
g1132 not 6442(1006) ; 6446(1332)
g1133 and 4175(1007) ; 6439(1333)
g1134 and 4175(1007) ; 7585(1334)
g1135 and 4172(1008) ; 6447(1335)
g1136 and 4172(1008) ; 7588(1336)
g1137 and 4169(1009) ; 6455(1337)
g1138 and 4169(1009) ; 7575(1338)
g1139 and 4157(1010) ; 6479(1339)
g1140 and 4157(1010) ; 7559(1340)
g1141 not 7554(1011) ; 7558(1341)
g1142 and 4511(1012) ; 7541(1342)
g1143 and 4511(1012) ; 7361(1343)
g1144 and 4508(1013) ; 7369(1344)
g1145 and 4508(1013) ; 7544(1345)
g1146 and 4505(1014) ; 7531(1346)
g1147 and 4505(1014) ; 7377(1347)
g1148 and 4502(1015) ; 7534(1348)
g1149 and 4502(1015) ; 7417(1349)
g1150 and 3833(1016) ; 6578(1350)
g1151 and 3833(1016) ; 6758(1351)
g1152 and 3833(1016) ; 6864(1352)
g1153 and 3810(823) 4172(1008) ; 3068(1353)
g1154 not 6450(1017) ; 6454(1354)
g1155 not 7242(1018) ; 7246(1355)
g1156 and 3801(824) 4163(994) ; 3090(1356)
g1157 not 6466(1019) ; 6470(1357)
g1158 not 7221(1020) ; 7227(1358)
g1159 and 3816(1021) ; 6602(1359)
g1160 and 3816(1021) ; 6737(1360)
g1161 and 3816(1021) ; 6880(1361)
g1162 or 7256(1022)* 7249(1024)* ; 4202(1362)
g1163 not 6768(1023) ; 6772(1363)
g1164 not 7249(1024) ; 7255(1364)
g1165 and 2320(1025) ; 6765(1365)
g1166 and 3173(717) 3170(866) ; 3222(1366)
g1167 or 3211(827)* 3210(1026)* ; 3212(1367)
g1168 or 5245(830)* 5242(917)* ; 1156(1368)
g1169 or 5237(720)* 5234(918)* ; 1152(1369)
g1170 and 3804(833) 4166(995) ; 3079(1370)
g1171 not 6498(1032) ; 6502(1371)
g1172 not 7232(1033) ; 7236(1372)
g1173 and 3821(1034) ; 6748(1373)
g1174 and 3821(1034) ; 6912(1374)
g1175 and 3821(1034) ; 6594(1375)
g1176 and 3828(1035) ; 6745(1376)
g1177 and 3828(1035) ; 6872(1377)
g1178 and 3828(1035) ; 6586(1378)
g1179 and 3807(834) 4169(1009) ; 3076(1379)
g1180 not 6458(1036) ; 6462(1380)
g1181 not 7229(1037) ; 7235(1381)
g1182 and 2323(1038) ; 5924(1382)
g1183 and 2323(1038) ; 6036(1383)
g1184 and 2323(1038) ; 6776(1384)
g1185 and 2308(835) 4490(1000) ; 4348(1385)
g1186 not 7412(1039) ; 7416(1386)
g1187 not 7260(1040) ; 7264(1387)
g1188 and 2329(1041) ; 6773(1388)
g1189 and 2329(1041) ; 6028(1389)
g1190 and 2329(1041) ; 5916(1390)
g1191 not 7404(1042) ; 7408(1391)
g1192 and 2312(836) 4493(998) ; 4341(1392)
g1193 not 7257(1043) ; 7263(1393)
g1194 and 2335(1044) ; 5908(1394)
g1195 and 2335(1044) ; 6020(1395)
g1196 and 2335(1044) ; 6784(1396)
g1197 and 2316(837) 4496(999) ; 4333(1397)
g1198 not 7396(1045) ; 7400(1398)
g1199 not 7268(1046) ; 7272(1399)
g1200 and 3695(1050) 3686(838) ; 4349(1400)
g1201 not 7425(1047) ; 7431(1401)
g1202 not 5929(1048) ; 5935(1402)
g1203 not 6049(1049) ; 6055(1403)
g1204 and 3695(1050) ; 7428(1404)
g1205 and 1535(302) 2320(1025) ; 4389(1405)
g1206 not 5284(1051) ; 5288(1406)
g1207 not 5300(1052) ; 5304(1407)
g1208 not 6530(1053) ; 6534(1408)
g1209 not 5289(1054) ; 5295(1409)
g1210 not 6538(1055) ; 6542(1410)
g1211 not 5292(1056) ; 5296(1411)
g1212 not 6546(1057) ; 6550(1412)
g1213 not 5281(1058) ; 5287(1413)
g1214 not 6562(1059) ; 6566(1414)
g1215 or 5312(1061)* 5305(845)* ; 5314(1415)
g1216 or 5311(1060)* 5308(846)* ; 5313(1416)
g1217 not 5297(1062) ; 5303(1417)
g1218 not 6522(1063) ; 6526(1418)
g1219 not 7327(1064) ; 7333(1419)
g1220 not 6370(1065) ; 6374(1420)
g1221 not 6378(1066) ; 6382(1421)
g1222 not 7330(1067) ; 7334(1422)
g1223 not 7317(1068) ; 7323(1423)
g1224 not 6386(1069) ; 6390(1424)
g1225 not 6426(1070) ; 6430(1425)
g1226 not 7320(1071) ; 7324(1426)
g1227 not 7309(1072) ; 7315(1427)
g1228 not 6394(1073) ; 6398(1428)
g1229 not 5339(1074) ; 5345(1429)
g1230 not 5764(1075) ; 5768(1430)
g1231 not 5412(1076) ; 5416(1431)
g1232 not 5452(1077) ; 5456(1432)
g1233 not 5772(1078) ; 5776(1433)
g1234 not 5342(1079) ; 5346(1434)
g1235 not 5331(1080) ; 5337(1435)
g1236 not 5780(1081) ; 5784(1436)
g1237 not 5420(1082) ; 5424(1437)
g1238 not 5349(1083) ; 5355(1438)
g1239 not 5396(1084) ; 5400(1439)
g1240 not 5748(1085) ; 5752(1440)
g1241 not 5756(1086) ; 5760(1441)
g1242 not 5404(1087) ; 5408(1442)
g1243 not 5352(1088) ; 5356(1443)
g1244 not 5202(1089) ; 5206(1444)
g1245 not 4892(1090) ; 4896(1445)
g1246 not 5266(1091) ; 5270(1446)
g1247 not 5255(1092) ; 5261(1447)
g1248 not 4900(1093) ; 4904(1448)
g1249 not 5210(1094) ; 5214(1449)
g1250 not 5218(1095) ; 5222(1450)
g1251 not 4908(1096) ; 4912(1451)
g1252 not 5258(1097) ; 5262(1452)
g1253 not 5247(1098) ; 5253(1453)
g1254 not 4924(1099) ; 4928(1454)
g1255 not 5226(1100) ; 5230(1455)
g1256 not 5250(1101) ; 5254(1456)
g1257 or 5278(1103)* 5271(863)* ; 5280(1457)
g1258 or 5277(1102)* 5274(864)* ; 5279(1458)
g1259 not 5263(1104) ; 5269(1459)
g1260 not 4884(1105) ; 4888(1460)
g1261 not 5194(1106) ; 5198(1461)
g1262 and 3170(866) 3212(1367) ; 3216(1462)
g1263 or 6859(431)* 6856(1327)* ; 3843(1463)
g1264 or 6573(432)* 6570(1329)* ; 3281(1464)
g1265 or 6581(433)* 6578(1350)* ; 3293(1465)
g1266 or 6867(434)* 6864(1352)* ; 3854(1466)
g1267 or 6589(435)* 6586(1378)* ; 3312(1467)
g1268 or 6875(436)* 6872(1377)* ; 3872(1468)
g1269 and 3335(1113) ; 6679(1469)
g1270 and 3891(1114) ; 6983(1470)
g1271 not 6925(1115) ; 6931(1471)
g1272 or 6915(437)* 6912(1374)* ; 3987(1472)
g1273 or 6597(438)* 6594(1375)* ; 3342(1473)
g1274 not 6671(1116) ; 6677(1474)
g1275 or 6883(439)* 6880(1361)* ; 3897(1475)
g1276 or 6605(440)* 6602(1359)* ; 3351(1476)
g1277 or 6613(441)* 6610(1266)* ; 3363(1477)
g1278 or 6891(442)* 6888(1267)* ; 3909(1478)
g1279 or 6899(443)* 6896(1302)* ; 3930(1479)
g1280 or 6621(444)* 6618(1303)* ; 3379(1480)
g1281 or 6907(445)* 6904(1296)* ; 3955(1481)
g1282 or 6629(446)* 6626(1297)* ; 3397(1482)
g1283 and 3979(1126) ; 7129(1483)
g1284 or 6637(447)* 6634(1275)* ; 3415(1484)
g1285 not 7041(1127) ; 7047(1485)
g1286 or 6923(448)* 6920(1276)* ; 3995(1486)
g1287 or 5991(449)* 5988(1290)* ; 2587(1487)
g1288 or 5871(450)* 5868(1291)* ; 2341(1488)
g1289 or 5879(451)* 5876(1259)* ; 2352(1489)
g1290 or 5999(452)* 5996(1260)* ; 2598(1490)
g1291 or 6007(453)* 6004(1254)* ; 2616(1491)
g1292 or 5887(454)* 5884(1255)* ; 2370(1492)
g1293 and 2391(1134) ; 5977(1493)
g1294 and 2635(1135) ; 6115(1494)
g1295 not 6057(1136) ; 6063(1495)
g1296 or 6047(455)* 6044(1251)* ; 2732(1496)
g1297 or 5895(456)* 5892(1250)* ; 2398(1497)
g1298 not 5969(1137) ; 5975(1498)
g1299 or 5903(457)* 5900(1288)* ; 2407(1499)
g1300 or 6015(458)* 6012(1287)* ; 2641(1500)
g1301 or 6023(459)* 6020(1395)* ; 2653(1501)
g1302 or 5911(460)* 5908(1394)* ; 2418(1502)
g1303 or 5919(461)* 5916(1390)* ; 2434(1503)
g1304 or 6031(462)* 6028(1389)* ; 2674(1504)
g1305 or 6039(463)* 6036(1383)* ; 2699(1505)
g1306 or 5927(464)* 5924(1382)* ; 2452(1506)
g1307 or 7504(1150)* 7497(868)* ; 7506(1507)
g1308 or 6374(1420)* 6367(869)* ; 2955(1508)
g1309 or 5400(1439)* 5393(352)* ; 1545(1509)
g1310 or 5752(1440)* 5745(353)* ; 1794(1510)
g1311 or 7503(1146)* 7500(873)* ; 7505(1511)
g1312 or 6382(1421)* 6375(874)* ; 2964(1512)
g1313 or 5760(1441)* 5753(354)* ; 1804(1513)
g1314 or 5408(1442)* 5401(355)* ; 1555(1514)
g1315 or 6390(1424)* 6383(880)* ; 2972(1515)
g1316 or 7494(1164)* 7487(881)* ; 7496(1516)
g1317 or 5416(1431)* 5409(356)* ; 1572(1517)
g1318 or 5768(1430)* 5761(357)* ; 1821(1518)
g1319 not 5523(1158) ; 5529(1519)
g1320 not 5857(1159) ; 5863(1520)
g1321 or 5776(1433)* 5769(358)* ; 1849(1521)
g1322 or 5456(1432)* 5449(359)* ; 1686(1522)
g1323 or 7493(1155)* 7490(887)* ; 7495(1523)
g1324 or 6430(1425)* 6423(888)* ; 3017(1524)
g1325 or 7486(1173)* 7479(890)* ; 4548(1525)
g1326 or 6398(1428)* 6391(891)* ; 2981(1526)
g1327 or 5424(1437)* 5417(360)* ; 1597(1527)
g1328 or 5784(1436)* 5777(361)* ; 1858(1528)
g1329 or 5792(1243)* 5785(362)* ; 1868(1529)
g1330 or 5432(1242)* 5425(363)* ; 1608(1530)
g1331 or 6406(1230)* 6399(897)* ; 2991(1531)
g1332 or 7485(1166)* 7482(898)* ; 4547(1532)
g1333 or 7478(1181)* 7471(902)* ; 4539(1533)
g1334 or 6414(1229)* 6407(903)* ; 3000(1534)
g1335 or 5440(1240)* 5433(364)* ; 1629(1535)
g1336 or 5800(1239)* 5793(365)* ; 1884(1536)
g1337 or 5808(1237)* 5801(366)* ; 1902(1537)
g1338 or 5448(1236)* 5441(367)* ; 1654(1538)
g1339 or 6422(1226)* 6415(907)* ; 3008(1539)
g1340 or 7477(1174)* 7474(908)* ; 4538(1540)
g1341 not 5669(1182) ; 5675(1541)
g1342 or 5464(1246)* 5457(368)* ; 1694(1542)
g1343 or 6438(1233)* 6431(914)* ; 3020(1543)
g1344 or 5816(1245)* 5809(369)* ; 1920(1544)
g1345 or 7469(1186)* 7466(771)* ; 4529(1545)
g1346 or 6720(1189)* 6719(1202)* ; 6832(1546)
g1347 or 953(1197) 917(1190) ; 4932(1547)
g1348 not 917(1190) ; 4973(1548)
g1349 not 4983(1191) ; 4987(1549)
g1350 not 908(1192) ; 912(1550)
g1351 or 914(1200) 913(1027) 777(370) ; 4942(1551)
g1352 not 1117(1193) ; 1121(1552)
g1353 not 1108(1196) ; 1112(1553)
g1354 not 902(1199) ; 906(1554)
g1355 not 4993(1203) ; 4997(1555)
g1356 not 4952(1204) ; 4956(1556)
g1357 or 6710(1213)* 6703(927)* ; 3521(1557)
g1358 or 6526(1418)* 6519(928)* ; 3175(1558)
g1359 or 4888(1460)* 4881(375)* ; 791(1559)
g1360 or 5198(1461)* 5191(376)* ; 1025(1560)
g1361 or 5206(1444)* 5199(377)* ; 1037(1561)
g1362 or 4896(1445)* 4889(378)* ; 804(1562)
g1363 or 6534(1408)* 6527(932)* ; 3185(1563)
g1364 or 6709(1206)* 6706(933)* ; 3520(1564)
g1365 or 5222(1450)* 5215(379)* ; 1073(1565)
g1366 or 6550(1412)* 6543(937)* ; 3202(1566)
g1367 or 6701(1281)* 6698(938)* ; 3511(1567)
g1368 or 4912(1451)* 4905(380)* ; 852(1568)
g1369 not 5099(1218) ; 5105(1569)
g1370 or 4928(1454)* 4921(381)* ; 894(1570)
g1371 or 6566(1414)* 6559(944)* ; 3214(1571)
g1372 or 5230(1455)* 5223(382)* ; 1092(1572)
g1373 or 6693(1222)* 6690(780)* ; 3502(1573)
g1374 or 7299(1232)* 7296(811)* ; 4224(1574)
g1375 or 6421(1180)* 6418(947)* ; 3007(1575)
g1376 or 7307(1228)* 7304(948)* ; 4233(1576)
g1377 or 7308(1227)* 7301(949)* ; 4234(1577)
g1378 or 6413(1175)* 6410(950)* ; 2999(1578)
g1379 or 6405(1172)* 6402(951)* ; 2990(1579)
g1380 or 7315(1427)* 7312(952)* ; 4242(1580)
g1381 or 6437(1187)* 6434(954)* ; 3019(1581)
g1382 or 5321(1244)* 5318(816)* ; 1261(1582)
g1383 or 5329(1238)* 5326(956)* ; 1270(1583)
g1384 or 5330(1235)* 5323(959)* ; 1271(1584)
g1385 or 5337(1435)* 5334(962)* ; 1279(1585)
g1386 not 7276(1247) ; 7280(1586)
g1387 not 7420(1249) ; 7424(1587)
g1388 not 5892(1250) ; 5896(1588)
g1389 not 6044(1251) ; 6048(1589)
g1390 not 6792(1252) ; 6796(1590)
g1391 not 6789(1253) ; 6795(1591)
g1392 not 6004(1254) ; 6008(1592)
g1393 not 5884(1255) ; 5888(1593)
g1394 not 7380(1257) ; 7384(1594)
g1395 not 7273(1258) ; 7279(1595)
g1396 not 5876(1259) ; 5880(1596)
g1397 not 5996(1260) ; 6000(1597)
g1398 not 6802(1261) ; 6806(1598)
g1399 not 7372(1263) ; 7376(1599)
g1400 not 7286(1264) ; 7290(1600)
g1401 not 6740(1265) ; 6744(1601)
g1402 not 6610(1266) ; 6614(1602)
g1403 not 6888(1267) ; 6892(1603)
g1404 not 6474(1269) ; 6478(1604)
g1405 or 7227(1358)* 7224(1270)* ; 4196(1605)
g1406 not 7224(1270) ; 7228(1606)
g1407 not 6506(1272) ; 6510(1607)
g1408 or 7212(1277)* 7205(1273)* ; 4179(1608)
g1409 not 7205(1273) ; 7211(1609)
g1410 or 6728(1278)* 6721(1274)* ; 3526(1610)
g1411 not 6721(1274) ; 6727(1611)
g1412 not 6634(1275) ; 6638(1612)
g1413 not 6920(1276) ; 6924(1613)
g1414 or 4904(1448)* 4897(548)* ; 826(1614)
g1415 or 5214(1449)* 5207(549)* ; 1054(1615)
g1416 or 6702(1216)* 6695(983)* ; 3512(1616)
g1417 or 6542(1410)* 6535(984)* ; 3194(1617)
g1418 not 7388(1283) ; 7392(1618)
g1419 or 7272(1399)* 7265(1285)* ; 4220(1619)
g1420 not 7265(1285) ; 7271(1620)
g1421 not 6781(1286) ; 6787(1621)
g1422 not 6012(1287) ; 6016(1622)
g1423 not 5900(1288) ; 5904(1623)
g1424 not 6799(1289) ; 6805(1624)
g1425 not 5988(1290) ; 5992(1625)
g1426 not 5868(1291) ; 5872(1626)
g1427 not 7364(1292) ; 7368(1627)
g1428 not 7283(1294) ; 7289(1628)
g1429 not 6732(1295) ; 6736(1629)
g1430 not 6904(1296) ; 6908(1630)
g1431 not 6626(1297) ; 6630(1631)
g1432 not 6490(1299) ; 6494(1632)
g1433 not 7216(1300) ; 7220(1633)
g1434 not 6729(1301) ; 6735(1634)
g1435 not 6896(1302) ; 6900(1635)
g1436 not 6618(1303) ; 6622(1636)
g1437 not 6482(1304) ; 6486(1637)
g1438 not 7213(1306) ; 7219(1638)
g1439 not 6471(1307) ; 6477(1639)
g1440 not 7570(1308) ; 7574(1640)
g1441 or 6470(1357)* 6463(1309)* ; 3081(1641)
g1442 not 6463(1309) ; 6469(1642)
g1443 not 7567(1310) ; 7573(1643)
g1444 or 6502(1371)* 6495(1311)* ; 3118(1644)
g1445 not 6495(1311) ; 6501(1645)
g1446 not 7578(1312) ; 7582(1646)
g1447 not 6487(1313) ; 6493(1647)
g1448 not 7562(1314) ; 7566(1648)
g1449 not 6503(1315) ; 6509(1649)
g1450 or 7558(1341)* 7551(1316)* ; 4576(1650)
g1451 not 7551(1316) ; 7557(1651)
g1452 not 7515(1317) ; 7521(1652)
g1453 or 7408(1391)* 7401(1318)* ; 4335(1653)
g1454 not 7401(1318) ; 7407(1654)
g1455 or 7400(1398)* 7393(1319)* ; 4326(1655)
g1456 not 7393(1319) ; 7399(1656)
g1457 not 7526(1320) ; 7530(1657)
g1458 or 7416(1386)* 7409(1321)* ; 4343(1658)
g1459 not 7409(1321) ; 7415(1659)
g1460 not 7518(1322) ; 7522(1660)
g1461 not 7523(1323) ; 7529(1661)
g1462 not 7385(1324) ; 7391(1662)
g1463 or 7514(1326)* 7507(1002)* ; 4553(1663)
g1464 or 7513(1325)* 7510(1003)* ; 4552(1664)
g1465 not 6856(1327) ; 6860(1665)
g1466 not 6755(1328) ; 6761(1666)
g1467 not 6570(1329) ; 6574(1667)
g1468 or 7246(1355)* 7239(1005)* ; 7248(1668)
g1469 or 6446(1332)* 6439(1333)* ; 3051(1669)
g1470 not 6439(1333) ; 6445(1670)
g1471 not 7585(1334) ; 7591(1671)
g1472 or 6454(1354)* 6447(1335)* ; 3061(1672)
g1473 not 6447(1335) ; 6453(1673)
g1474 not 7588(1336) ; 7592(1674)
g1475 or 6462(1380)* 6455(1337)* ; 3070(1675)
g1476 not 6455(1337) ; 6461(1676)
g1477 not 7575(1338) ; 7581(1677)
g1478 not 6479(1339) ; 6485(1678)
g1479 not 7559(1340) ; 7565(1679)
g1480 not 7541(1342) ; 7547(1680)
g1481 not 7361(1343) ; 7367(1681)
g1482 not 7369(1344) ; 7375(1682)
g1483 not 7544(1345) ; 7548(1683)
g1484 not 7531(1346) ; 7537(1684)
g1485 not 7377(1347) ; 7383(1685)
g1486 not 7534(1348) ; 7538(1686)
g1487 not 7417(1349) ; 7423(1687)
g1488 not 6578(1350) ; 6582(1688)
g1489 not 6758(1351) ; 6762(1689)
g1490 not 6864(1352) ; 6868(1690)
g1491 or 7245(1331)* 7242(1018)* ; 7247(1691)
g1492 not 6602(1359) ; 6606(1692)
g1493 not 6737(1360) ; 6743(1693)
g1494 not 6880(1361) ; 6884(1694)
g1495 or 7255(1364)* 7252(825)* ; 4201(1695)
g1496 or 6772(1363)* 6765(1365)* ; 3549(1696)
g1497 not 6765(1365) ; 6771(1697)
g1498 or 3222(1366) 3221(557) ; 3223(1698)
g1499 or 5246(1194)* 5239(719)* ; 1157(1699)
g1500 or 5238(1195)* 5231(561)* ; 1153(1700)
g1501 or 7235(1381)* 7232(1033)* ; 7237(1701)
g1502 not 6748(1373) ; 6752(1702)
g1503 not 6912(1374) ; 6916(1703)
g1504 not 6594(1375) ; 6598(1704)
g1505 not 6745(1376) ; 6751(1705)
g1506 not 6872(1377) ; 6876(1706)
g1507 not 6586(1378) ; 6590(1707)
g1508 or 7236(1372)* 7229(1037)* ; 7238(1708)
g1509 not 5924(1382) ; 5928(1709)
g1510 not 6036(1383) ; 6040(1710)
g1511 not 6776(1384) ; 6780(1711)
g1512 or 7263(1393)* 7260(1040)* ; 4210(1712)
g1513 not 6773(1388) ; 6779(1713)
g1514 not 6028(1389) ; 6032(1714)
g1515 not 5916(1390) ; 5920(1715)
g1516 or 7264(1387)* 7257(1043)* ; 4211(1716)
g1517 not 5908(1394) ; 5912(1717)
g1518 not 6020(1395) ; 6024(1718)
g1519 not 6784(1396) ; 6788(1719)
g1520 or 7431(1401)* 7428(1404)* ; 4353(1720)
g1521 and 4389(1405) 3682(839) ; 2481(1721)
g1522 and 4389(1405) 3682(839) ; 2724(1722)
g1523 and 4389(1405)* 3682(839)* ; 6173(1723)
g1524 not 7428(1404) ; 7432(1724)
g1525 and 4389(1405) ; 6052(1725)
g1526 and 4389(1405) ; 5932(1726)
g1527 or 5287(1413)* 5284(1051)* ; 1238(1727)
g1528 or 5303(1417)* 5300(1052)* ; 1256(1728)
g1529 or 6533(1212)* 6530(1053)* ; 3184(1729)
g1530 or 5296(1411)* 5289(1054)* ; 1248(1730)
g1531 or 6541(1282)* 6538(1055)* ; 3193(1731)
g1532 or 5295(1409)* 5292(1056)* ; 1247(1732)
g1533 or 6549(1215)* 6546(1057)* ; 3201(1733)
g1534 or 5288(1406)* 5281(1058)* ; 1239(1734)
g1535 or 6565(1223)* 6562(1059)* ; 3213(1735)
g1536 or 5314(1415)* 5313(1416)* ; 5380(1736)
g1537 or 5304(1407)* 5297(1062)* ; 1257(1737)
g1538 or 6525(1207)* 6522(1063)* ; 3174(1738)
g1539 or 7334(1422)* 7327(1064)* ; 7336(1739)
g1540 or 6373(1147)* 6370(1065)* ; 2954(1740)
g1541 or 6381(1151)* 6378(1066)* ; 2963(1741)
g1542 or 7333(1419)* 7330(1067)* ; 7335(1742)
g1543 or 7324(1426)* 7317(1068)* ; 7326(1743)
g1544 or 6389(1154)* 6386(1069)* ; 2971(1744)
g1545 or 6429(1165)* 6426(1070)* ; 3016(1745)
g1546 or 7323(1423)* 7320(1071)* ; 7325(1746)
g1547 or 7316(1231)* 7309(1072)* ; 4243(1747)
g1548 or 6397(1167)* 6394(1073)* ; 2980(1748)
g1549 or 5346(1434)* 5339(1074)* ; 5348(1749)
g1550 or 5345(1429)* 5342(1079)* ; 5347(1750)
g1551 or 5338(1241)* 5331(1080)* ; 1280(1751)
g1552 or 5356(1443)* 5349(1083)* ; 5358(1752)
g1553 or 5355(1438)* 5352(1088)* ; 5357(1753)
g1554 or 5269(1459)* 5266(1091)* ; 1233(1754)
g1555 or 5262(1452)* 5255(1092)* ; 1225(1755)
g1556 or 5261(1447)* 5258(1097)* ; 1224(1756)
g1557 or 5254(1456)* 5247(1098)* ; 1216(1757)
g1558 or 5253(1453)* 5250(1101)* ; 1215(1758)
g1559 or 5280(1457)* 5279(1458)* ; 5372(1759)
g1560 or 5270(1446)* 5263(1104)* ; 1234(1760)
g1561 not 3216(1462) ; 3220(1761)
g1562 or 6860(1665)* 6853(318)* ; 3844(1762)
g1563 or 6574(1667)* 6567(319)* ; 3282(1763)
g1564 or 6582(1688)* 6575(320)* ; 3294(1764)
g1565 or 6868(1690)* 6861(321)* ; 3855(1765)
g1566 or 6590(1707)* 6583(322)* ; 3313(1766)
g1567 or 6876(1706)* 6869(323)* ; 3873(1767)
g1568 not 6679(1469) ; 6685(1768)
g1569 not 6983(1470) ; 6989(1769)
g1570 or 6916(1703)* 6909(324)* ; 3988(1770)
g1571 or 6598(1704)* 6591(325)* ; 3343(1771)
g1572 or 6884(1694)* 6877(326)* ; 3898(1772)
g1573 or 6606(1692)* 6599(327)* ; 3352(1773)
g1574 or 6614(1602)* 6607(328)* ; 3364(1774)
g1575 or 6892(1603)* 6885(329)* ; 3910(1775)
g1576 or 6900(1635)* 6893(330)* ; 3931(1776)
g1577 or 6622(1636)* 6615(331)* ; 3380(1777)
g1578 or 6908(1630)* 6901(332)* ; 3956(1778)
g1579 or 6630(1631)* 6623(333)* ; 3398(1779)
g1580 not 7129(1483) ; 7135(1780)
g1581 or 6638(1612)* 6631(334)* ; 3416(1781)
g1582 or 6924(1613)* 6917(335)* ; 3996(1782)
g1583 or 5992(1625)* 5985(336)* ; 2588(1783)
g1584 or 5872(1626)* 5865(337)* ; 2342(1784)
g1585 or 5880(1596)* 5873(338)* ; 2353(1785)
g1586 or 6000(1597)* 5993(339)* ; 2599(1786)
g1587 or 6008(1592)* 6001(340)* ; 2617(1787)
g1588 or 5888(1593)* 5881(341)* ; 2371(1788)
g1589 not 5977(1493) ; 5983(1789)
g1590 not 6115(1494) ; 6121(1790)
g1591 or 6048(1589)* 6041(342)* ; 2733(1791)
g1592 or 5896(1588)* 5889(343)* ; 2399(1792)
g1593 or 5904(1623)* 5897(344)* ; 2408(1793)
g1594 or 6016(1622)* 6009(345)* ; 2642(1794)
g1595 or 6024(1718)* 6017(346)* ; 2654(1795)
g1596 or 5912(1717)* 5905(347)* ; 2419(1796)
g1597 or 5920(1715)* 5913(348)* ; 2435(1797)
g1598 or 6032(1714)* 6025(349)* ; 2675(1798)
g1599 or 6040(1710)* 6033(350)* ; 2700(1799)
g1600 or 5928(1709)* 5921(351)* ; 2453(1800)
g1601 or 7506(1507)* 7505(1511)* ; 7595(1801)
g1602 or 2955(1508)* 2954(1740)* ; 2956(1802)
g1603 or 1545(1509)* 1544(1148)* ; 1546(1803)
g1604 or 1794(1510)* 1793(1149)* ; 1795(1804)
g1605 or 2964(1512)* 2963(1741)* ; 2965(1805)
g1606 or 1804(1513)* 1803(1152)* ; 1805(1806)
g1607 or 1555(1514)* 1554(1153)* ; 1556(1807)
g1608 or 2972(1515)* 2971(1744)* ; 2973(1808)
g1609 or 7496(1516)* 7495(1523)* ; 7598(1809)
g1610 or 1572(1517)* 1571(1156)* ; 1573(1810)
g1611 or 1821(1518)* 1820(1157)* ; 1822(1811)
g1612 or 1849(1521)* 1848(1160)* ; 1850(1812)
g1613 or 1686(1522)* 1685(1163)* ; 1687(1813)
g1614 or 3017(1524)* 3016(1745)* ; 3018(1814)
g1615 or 4548(1525)* 4547(1532)* ; 4549(1815)
g1616 or 2981(1526)* 2980(1748)* ; 2982(1816)
g1617 or 1597(1527)* 1596(1168)* ; 1598(1817)
g1618 or 1858(1528)* 1857(1169)* ; 1859(1818)
g1619 or 1868(1529)* 1867(1170)* ; 1869(1819)
g1620 or 1608(1530)* 1607(1171)* ; 1609(1820)
g1621 or 2991(1531)* 2990(1579)* ; 2992(1821)
g1622 or 4539(1533)* 4538(1540)* ; 4540(1822)
g1623 or 3000(1534)* 2999(1578)* ; 3001(1823)
g1624 or 1629(1535)* 1628(1176)* ; 1630(1824)
g1625 or 1884(1536)* 1883(1177)* ; 1885(1825)
g1626 or 1902(1537)* 1901(1178)* ; 1903(1826)
g1627 or 1654(1538)* 1653(1179)* ; 1655(1827)
g1628 or 3008(1539)* 3007(1575)* ; 3009(1828)
g1629 or 1694(1542)* 1693(1184)* ; 1695(1829)
g1630 or 4530(1185)* 4529(1545)* ; 4531(1830)
g1631 or 3020(1543)* 3019(1581)* ; 3021(1831)
g1632 or 1920(1544)* 1919(1188)* ; 1921(1832)
g1633 not 6832(1546) ; 6836(1833)
g1634 not 4932(1547) ; 4936(1834)
g1635 not 4973(1548) ; 4977(1835)
g1636 or 906(1554)* 912(1550)* ; 957(1836)
g1637 not 4942(1551) ; 4946(1837)
g1638 or 1112(1553)* 1121(1552)* ; 1176(1838)
g1639 or 3521(1557)* 3520(1564)* ; 3522(1839)
g1640 or 3175(1558)* 3174(1738)* ; 3176(1840)
g1641 or 791(1559)* 790(1208)* ; 792(1841)
g1642 or 1025(1560)* 1024(1209)* ; 1026(1842)
g1643 or 1037(1561)* 1036(1210)* ; 1038(1843)
g1644 or 804(1562)* 803(1211)* ; 805(1844)
g1645 or 3185(1563)* 3184(1729)* ; 3186(1845)
g1646 or 1073(1565)* 1072(1214)* ; 1074(1846)
g1647 or 3202(1566)* 3201(1733)* ; 3203(1847)
g1648 or 3512(1616)* 3511(1567)* ; 3513(1848)
g1649 or 852(1568)* 851(1217)* ; 853(1849)
g1650 or 894(1570)* 893(1220)* ; 895(1850)
g1651 or 3503(1221)* 3502(1573)* ; 3504(1851)
g1652 or 3214(1571)* 3213(1735)* ; 3215(1852)
g1653 or 1092(1572)* 1091(1224)* ; 1093(1853)
g1654 or 4225(1225)* 4224(1574)* ; 4226(1854)
g1655 or 4234(1577)* 4233(1576)* ; 4235(1855)
g1656 or 4243(1747)* 4242(1580)* ; 4244(1856)
g1657 or 1262(1234)* 1261(1582)* ; 1263(1857)
g1658 or 1271(1584)* 1270(1583)* ; 1272(1858)
g1659 or 1280(1751)* 1279(1585)* ; 1281(1859)
g1660 or 7279(1595)* 7276(1247)* ; 7281(1860)
g1661 or 7423(1687)* 7420(1249)* ; 4350(1861)
g1662 or 6795(1591)* 6792(1252)* ; 6797(1862)
g1663 or 6796(1590)* 6789(1253)* ; 6798(1863)
g1664 or 7383(1685)* 7380(1257)* ; 4306(1864)
g1665 or 7280(1586)* 7273(1258)* ; 7282(1865)
g1666 or 6805(1624)* 6802(1261)* ; 6807(1866)
g1667 or 7375(1682)* 7372(1263)* ; 4298(1867)
g1668 or 7289(1628)* 7286(1264)* ; 7291(1868)
g1669 or 6743(1693)* 6740(1265)* ; 3543(1869)
g1670 or 6477(1639)* 6474(1269)* ; 3091(1870)
g1671 or 6509(1649)* 6506(1272)* ; 3120(1871)
g1672 or 7211(1609)* 7208(978)* ; 4178(1872)
g1673 or 6727(1611)* 6724(979)* ; 3525(1873)
g1674 or 826(1614)* 825(1279)* ; 827(1874)
g1675 or 1054(1615)* 1053(1280)* ; 1055(1875)
g1676 or 3194(1617)* 3193(1731)* ; 3195(1876)
g1677 or 7391(1662)* 7388(1283)* ; 4315(1877)
g1678 or 6788(1719)* 6781(1286)* ; 3567(1878)
g1679 or 6806(1598)* 6799(1289)* ; 6808(1879)
g1680 or 7367(1681)* 7364(1292)* ; 4289(1880)
g1681 or 7290(1600)* 7283(1294)* ; 7292(1881)
g1682 or 6735(1634)* 6732(1295)* ; 3534(1882)
g1683 or 6493(1647)* 6490(1299)* ; 3108(1883)
g1684 or 7219(1638)* 7216(1300)* ; 4187(1884)
g1685 or 6736(1629)* 6729(1301)* ; 3535(1885)
g1686 or 6485(1678)* 6482(1304)* ; 3100(1886)
g1687 or 7220(1633)* 7213(1306)* ; 4188(1887)
g1688 or 6478(1604)* 6471(1307)* ; 3092(1888)
g1689 or 7573(1643)* 7570(1308)* ; 4593(1889)
g1690 or 7574(1640)* 7567(1310)* ; 4594(1890)
g1691 or 7581(1677)* 7578(1312)* ; 7583(1891)
g1692 or 6494(1632)* 6487(1313)* ; 3109(1892)
g1693 or 7565(1679)* 7562(1314)* ; 4584(1893)
g1694 or 6510(1607)* 6503(1315)* ; 3121(1894)
g1695 or 7522(1660)* 7515(1317)* ; 4562(1895)
g1696 or 7529(1661)* 7526(1320)* ; 4570(1896)
g1697 or 7521(1652)* 7518(1322)* ; 4561(1897)
g1698 or 7530(1657)* 7523(1323)* ; 4571(1898)
g1699 or 7392(1618)* 7385(1324)* ; 4316(1899)
g1700 or 4553(1663)* 4552(1664)* ; 4554(1900)
g1701 or 6762(1689)* 6755(1328)* ; 6764(1901)
g1702 or 7248(1668)* 7247(1691)* ; 7337(1902)
g1703 or 6445(1670)* 6442(1006)* ; 3050(1903)
g1704 or 7592(1674)* 7585(1334)* ; 7594(1904)
g1705 or 7591(1671)* 7588(1336)* ; 7593(1905)
g1706 or 7582(1646)* 7575(1338)* ; 7584(1906)
g1707 or 6486(1637)* 6479(1339)* ; 3101(1907)
g1708 or 7566(1648)* 7559(1340)* ; 4585(1908)
g1709 or 7557(1651)* 7554(1011)* ; 4575(1909)
g1710 or 7548(1683)* 7541(1342)* ; 7550(1910)
g1711 or 7368(1627)* 7361(1343)* ; 4290(1911)
g1712 or 7376(1599)* 7369(1344)* ; 4299(1912)
g1713 or 7547(1680)* 7544(1345)* ; 7549(1913)
g1714 or 7538(1686)* 7531(1346)* ; 7540(1914)
g1715 or 7384(1594)* 7377(1347)* ; 4307(1915)
g1716 or 7537(1684)* 7534(1348)* ; 7539(1916)
g1717 or 7424(1587)* 7417(1349)* ; 4351(1917)
g1718 or 6761(1666)* 6758(1351)* ; 6763(1918)
g1719 or 6453(1673)* 6450(1017)* ; 3060(1919)
g1720 or 6469(1642)* 6466(1019)* ; 3080(1920)
g1721 or 7228(1606)* 7221(1020)* ; 4197(1921)
g1722 or 6744(1601)* 6737(1360)* ; 3544(1922)
g1723 or 4202(1362)* 4201(1695)* ; 4203(1923)
g1724 or 6771(1697)* 6768(1023)* ; 3548(1924)
g1725 not 3223(1698) ; 3227(1925)
g1726 or 4976(829)* 4973(1548)* ; 4978(1926)
g1727 or 1157(1699)* 1156(1368)* ; 1158(1927)
g1728 or 1153(1700)* 1152(1369)* ; 1154(1928)
g1729 or 4935(722)* 4932(1547)* ; 4937(1929)
g1730 or 6501(1645)* 6498(1032)* ; 3117(1930)
g1731 or 7238(1708)* 7237(1701)* ; 7340(1931)
g1732 or 6751(1705)* 6748(1373)* ; 6753(1932)
g1733 or 6752(1702)* 6745(1376)* ; 6754(1933)
g1734 or 6461(1676)* 6458(1036)* ; 3069(1934)
g1735 or 6779(1713)* 6776(1384)* ; 3557(1935)
g1736 or 7415(1659)* 7412(1039)* ; 4342(1936)
g1737 or 4211(1716)* 4210(1712)* ; 4212(1937)
g1738 or 6780(1711)* 6773(1388)* ; 3558(1938)
g1739 or 7407(1654)* 7404(1042)* ; 4334(1939)
g1740 or 6787(1621)* 6784(1396)* ; 3566(1940)
g1741 or 7399(1656)* 7396(1045)* ; 4325(1941)
g1742 or 7271(1620)* 7268(1046)* ; 4219(1942)
g1743 or 7432(1724)* 7425(1047)* ; 4354(1943)
g1744 and 2724(1722) ; 6261(1944)
g1745 or 5935(1402)* 5932(1726)* ; 2470(1945)
g1746 not 6173(1723) ; 6179(1946)
g1747 or 6055(1403)* 6052(1725)* ; 2740(1947)
g1748 not 6052(1725) ; 6056(1948)
g1749 not 5932(1726) ; 5936(1949)
g1750 or 1239(1734)* 1238(1727)* ; 1240(1950)
g1751 or 1257(1737)* 1256(1728)* ; 1258(1951)
g1752 or 1248(1730)* 1247(1732)* ; 1249(1952)
g1753 not 5380(1736) ; 5384(1953)
g1754 or 7336(1739)* 7335(1742)* ; 7353(1954)
g1755 or 7326(1743)* 7325(1746)* ; 7356(1955)
g1756 or 5348(1749)* 5347(1750)* ; 5362(1956)
g1757 or 5358(1752)* 5357(1753)* ; 5359(1957)
g1758 or 1234(1760)* 1233(1754)* ; 1235(1958)
g1759 or 1225(1755)* 1224(1756)* ; 1226(1959)
g1760 or 1216(1757)* 1215(1758)* ; 1217(1960)
g1761 not 5372(1759) ; 5376(1961)
g1762 or 3220(1761)* 3227(1925)* ; 3244(1962)
g1763 or 3844(1762)* 3843(1463)* ; 3845(1963)
g1764 or 3282(1763)* 3281(1464)* ; 3283(1964)
g1765 or 3294(1764)* 3293(1465)* ; 3295(1965)
g1766 or 3855(1765)* 3854(1466)* ; 3856(1966)
g1767 or 3313(1766)* 3312(1467)* ; 3314(1967)
g1768 or 3873(1767)* 3872(1468)* ; 3874(1968)
g1769 or 3988(1770)* 3987(1472)* ; 3989(1969)
g1770 or 3343(1771)* 3342(1473)* ; 3344(1970)
g1771 or 3898(1772)* 3897(1475)* ; 3899(1971)
g1772 or 3352(1773)* 3351(1476)* ; 3353(1972)
g1773 or 3364(1774)* 3363(1477)* ; 3365(1973)
g1774 or 3910(1775)* 3909(1478)* ; 3911(1974)
g1775 or 3931(1776)* 3930(1479)* ; 3932(1975)
g1776 or 3380(1777)* 3379(1480)* ; 3381(1976)
g1777 or 3956(1778)* 3955(1481)* ; 3957(1977)
g1778 or 3398(1779)* 3397(1482)* ; 3399(1978)
g1779 or 3416(1781)* 3415(1484)* ; 3417(1979)
g1780 or 3996(1782)* 3995(1486)* ; 3997(1980)
g1781 or 2588(1783)* 2587(1487)* ; 2589(1981)
g1782 or 2342(1784)* 2341(1488)* ; 2343(1982)
g1783 or 2353(1785)* 2352(1489)* ; 2354(1983)
g1784 or 2599(1786)* 2598(1490)* ; 2600(1984)
g1785 or 2617(1787)* 2616(1491)* ; 2618(1985)
g1786 or 2371(1788)* 2370(1492)* ; 2372(1986)
g1787 or 2733(1791)* 2732(1496)* ; 2734(1987)
g1788 or 2399(1792)* 2398(1497)* ; 2400(1988)
g1789 or 2408(1793)* 2407(1499)* ; 2409(1989)
g1790 or 2642(1794)* 2641(1500)* ; 2643(1990)
g1791 or 2654(1795)* 2653(1501)* ; 2655(1991)
g1792 or 2419(1796)* 2418(1502)* ; 2420(1992)
g1793 or 2435(1797)* 2434(1503)* ; 2436(1993)
g1794 or 2675(1798)* 2674(1504)* ; 2676(1994)
g1795 or 2700(1799)* 2699(1505)* ; 2701(1995)
g1796 or 2453(1800)* 2452(1506)* ; 2454(1996)
g1797 not 7595(1801) ; 7601(1997)
g1798 and 2956(1802) 2965(1805) 2973(1808) 3018(1814) ; 3022(1998)
g1799 and 1546(1803) 1556(1807) 1573(1810) 1687(1813) ; 1702(1999)
g1800 and 1546(1803) ; 5566(2000)
g1801 and 1546(1803) ; 5508(2001)
g1802 and 1795(1804) ; 5820(2002)
g1803 and 1795(1804) ; 5828(2003)
g1804 and 1795(1804) 1822(1811) 1850(1812) 1805(1806) ; 1935(2004)
g1805 and 2970(872) 2956(1802) ; 3025(2005)
g1806 and 1816(875) 1795(1804) ; 1938(2006)
g1807 and 1805(1806) ; 5844(2007)
g1808 and 1805(1806) ; 5836(2008)
g1809 and 1805(1806) 1822(1811) 1850(1812) ; 1944(2009)
g1810 and 1567(876) 1546(1803) ; 1705(2010)
g1811 and 1556(1807) ; 5518(2011)
g1812 and 1556(1807) 1573(1810) 1687(1813) ; 1711(2012)
g1813 and 1556(1807) ; 5576(2013)
g1814 and 1584(877) 1556(1807) ; 1712(2014)
g1815 and 1584(877) 1546(1803) 1556(1807) ; 1706(2015)
g1816 and 1584(877) 1556(1807) ; 1709(2016)
g1817 and 1834(878) 1795(1804) 1805(1806) ; 1939(2017)
g1818 and 1834(878) 1805(1806) ; 1942(2018)
g1819 and 1834(878) 1805(1806) ; 1945(2019)
g1820 and 2977(879) 2956(1802) 2965(1805) ; 3026(2020)
g1821 not 7598(1809) ; 7602(2021)
g1822 and 1573(1810) 1687(1813) ; 1749(2022)
g1823 and 1573(1810) ; 5498(2023)
g1824 and 1573(1810) ; 5556(2024)
g1825 and 1822(1811) ; 5860(2025)
g1826 and 1822(1811) ; 5852(2026)
g1827 and 1822(1811) 1850(1812) ; 1948(2027)
g1828 and 1556(1807) 1590(882) 1573(1810) ; 1710(2028)
g1829 and 1556(1807) 1590(882) 1546(1803) 1573(1810) ; 1707(2029)
g1830 and 1556(1807) 1590(882) 1573(1810) ; 1713(2030)
g1831 and 1590(882) 1573(1810) ; 1714(2031)
g1832 and 1805(1806) 1841(883) 1795(1804) 1822(1811) ; 1940(2032)
g1833 and 1805(1806) 1822(1811) 1841(883) ; 1946(2033)
g1834 and 1805(1806) 1841(883) 1822(1811) ; 1943(2034)
g1835 and 1841(883) 1822(1811) ; 1947(2035)
g1836 and 1841(883) 1822(1811) ; 1949(2036)
g1837 not 1850(1812) ; 1856(2037)
g1838 and 1687(1813) ; 5546(2038)
g1839 and 1687(1813) ; 5488(2039)
g1840 and 2965(1805) 2979(886) 2956(1802) 2973(1808) ; 3027(2040)
g1841 and 4549(1815) ; 4602(2041)
g1842 and 4549(1815) ; 4598(2042)
g1843 and 2982(1816) 2992(1821) 3001(1823) 3009(1828) 3021(1831) ; 3029(2043)
g1844 and 1598(1817) ; 5722(2044)
g1845 and 1598(1817) ; 5634(2045)
g1846 and 1598(1817) 1609(1820) 1630(1824) 1655(1827) 1695(1829) ; 1718(2046)
g1847 and 1903(1826) 1859(1818) 1885(1825) 1921(1832) 1869(1819) ; 1950(2047)
g1848 and 1859(1818) ; 4724(2048)
g1849 and 1624(894) 1598(1817) ; 1722(2049)
g1850 and 1880(895) 1859(1818) ; 1953(2050)
g1851 and 1869(1819) ; 4732(2051)
g1852 and 1609(1820) ; 5664(2052)
g1853 and 1655(1827) 1609(1820) 1630(1824) 1695(1829) ; 1736(2053)
g1854 and 1609(1820) ; 5654(2054)
g1855 and 2998(896) 2982(1816) ; 3030(2055)
g1856 and 1647(899) 1609(1820) ; 1737(2056)
g1857 and 1647(899) 1609(1820) ; 1733(2057)
g1858 and 1647(899) 1598(1817) 1609(1820) ; 1723(2058)
g1859 and 1897(900) 1869(1819) ; 1960(2059)
g1860 and 1897(900) 1859(1818) 1869(1819) ; 1954(2060)
g1861 and 3006(901) 2982(1816) 2992(1821) ; 3031(2061)
g1862 not 4540(1822) ; 4544(2062)
g1863 and 1630(1824) ; 5732(2063)
g1864 and 1630(1824) ; 5644(2064)
g1865 and 1655(1827) 1630(1824) 1695(1829) ; 1742(2065)
g1866 and 1885(1825) ; 4740(2066)
g1867 and 1609(1820) 1669(904) 1630(1824) ; 1738(2067)
g1868 and 1609(1820) 1669(904) 1630(1824) ; 1734(2068)
g1869 and 1609(1820) 1669(904) 1598(1817) 1630(1824) ; 1724(2069)
g1870 and 1669(904) 1630(1824) ; 1743(2070)
g1871 and 1669(904) 1630(1824) ; 1740(2071)
g1872 and 1869(1819) 1914(905) 1885(1825) ; 1961(2072)
g1873 and 1869(1819) 1914(905) 1859(1818) 1885(1825) ; 1955(2073)
g1874 and 1885(1825) 1914(905) ; 1965(2074)
g1875 and 1903(1826) ; 4748(2075)
g1876 and 1655(1827) ; 5624(2076)
g1877 and 1655(1827) ; 5712(2077)
g1878 and 1655(1827) 1695(1829) ; 1750(2078)
g1879 and 2992(1821) 3013(906) 2982(1816) 3001(1823) ; 3032(2079)
g1880 and 1609(1820) 1677(909) 1630(1824) 1655(1827) ; 1735(2080)
g1881 and 1609(1820) 1677(909) 1598(1817) 1630(1824) 1655(1827) ; 1725(2081)
g1882 and 1609(1820) 1677(909) 1630(1824) 1655(1827) ; 1739(2082)
g1883 and 1677(909) 1630(1824) 1655(1827) ; 1741(2083)
g1884 and 1677(909) 1655(1827) ; 1745(2084)
g1885 and 1677(909) 1630(1824) 1655(1827) ; 1744(2085)
g1886 and 1869(1819) 1929(910) 1885(1825) 1903(1826) ; 1962(2086)
g1887 and 1869(1819) 1929(910) 1859(1818) 1885(1825) 1903(1826) ; 1956(2087)
g1888 and 1929(910) 1903(1826) ; 1969(2088)
g1889 and 1929(910) 1885(1825) 1903(1826) ; 1966(2089)
g1890 and 1695(1829) ; 5702(2090)
g1891 and 1695(1829) ; 5614(2091)
g1892 and 2992(1821) 3015(912) 2982(1816) 3001(1823) 3009(1828) ; 3033(2092)
g1893 not 4531(1830) ; 4535(2093)
g1894 and 1921(1832) ; 4716(2094)
g1895 and 3522(1839) ; 3575(2095)
g1896 and 3522(1839) ; 3571(2096)
g1897 and 3176(1840) 3186(1845) 3195(1876) 3203(1847) 3215(1852) ; 3228(2097)
g1898 and 792(1841) ; 5152(2098)
g1899 and 792(1841) ; 5064(2099)
g1900 and 792(1841) 805(1844) 827(1874) 853(1849) 895(1850) ; 920(2100)
g1901 and 1074(1846) 1026(1842) 1055(1875) 1093(1853) 1038(1843) ; 1122(2101)
g1902 and 1026(1842) ; 4764(2102)
g1903 and 821(929) 792(1841) ; 925(2103)
g1904 and 1050(930) 1026(1842) ; 1125(2104)
g1905 and 1038(1843) ; 4772(2105)
g1906 and 805(1844) ; 5094(2106)
g1907 and 853(1849) 805(1844) 827(1874) 895(1850) ; 940(2107)
g1908 and 805(1844) ; 5084(2108)
g1909 and 3192(931) 3176(1840) ; 3231(2109)
g1910 and 805(1844) 868(934) 827(1874) ; 942(2110)
g1911 and 805(1844) 868(934) 827(1874) ; 938(2111)
g1912 and 805(1844) 868(934) 792(1841) 827(1874) ; 927(2112)
g1913 and 868(934) 827(1874) ; 947(2113)
g1914 and 868(934) 827(1874) ; 944(2114)
g1915 and 1038(1843) 1086(935) 1055(1875) ; 1133(2115)
g1916 and 1038(1843) 1086(935) 1026(1842) 1055(1875) ; 1127(2116)
g1917 and 1055(1875) 1086(935) ; 1137(2117)
g1918 and 1074(1846) ; 4788(2118)
g1919 and 3186(1845) 3207(936) 3176(1840) 3195(1876) ; 3233(2119)
g1920 not 3513(1848) ; 3517(2120)
g1921 and 853(1849) ; 5054(2121)
g1922 and 853(1849) 827(1874) 895(1850) ; 946(2122)
g1923 and 853(1849) ; 5142(2123)
g1924 and 853(1849) 895(1850) ; 956(2124)
g1925 and 805(1844) 877(939) 827(1874) 853(1849) ; 939(2125)
g1926 and 805(1844) 877(939) 792(1841) 827(1874) 853(1849) ; 928(2126)
g1927 and 805(1844) 877(939) 827(1874) 853(1849) ; 943(2127)
g1928 and 877(939) 827(1874) 853(1849) ; 945(2128)
g1929 and 877(939) 853(1849) ; 949(2129)
g1930 and 877(939) 827(1874) 853(1849) ; 948(2130)
g1931 and 1038(1843) 1102(940) 1055(1875) 1074(1846) ; 1134(2131)
g1932 and 1038(1843) 1102(940) 1026(1842) 1055(1875) 1074(1846) ; 1128(2132)
g1933 and 1102(940) 1074(1846) ; 1141(2133)
g1934 and 1102(940) 1055(1875) 1074(1846) ; 1138(2134)
g1935 and 895(1850) ; 5132(2135)
g1936 and 895(1850) ; 5044(2136)
g1937 and 3186(1845) 3209(942) 3176(1840) 3195(1876) 3203(1847) ; 3234(2137)
g1938 not 3504(1851) ; 3508(2138)
g1939 and 1093(1853) ; 4756(2139)
g1940 not 4226(1854) ; 4230(2140)
g1941 not 4235(1855) ; 4239(2141)
g1942 and 4244(1856) ; 4263(2142)
g1943 and 4244(1856) ; 4267(2143)
g1944 not 1263(1857) ; 1267(2144)
g1945 not 1272(1858) ; 1276(2145)
g1946 and 1281(1859) ; 1300(2146)
g1947 and 1281(1859) ; 1304(2147)
g1948 or 7282(1865)* 7281(1860)* ; 7348(2148)
g1949 or 4351(1917)* 4350(1861)* ; 4352(2149)
g1950 or 6798(1863)* 6797(1862)* ; 6822(2150)
g1951 or 4307(1915)* 4306(1864)* ; 4308(2151)
g1952 or 6808(1879)* 6807(1866)* ; 6819(2152)
g1953 or 4299(1912)* 4298(1867)* ; 4300(2153)
g1954 or 7292(1881)* 7291(1868)* ; 7345(2154)
g1955 or 3544(1922)* 3543(1869)* ; 3545(2155)
g1956 or 3092(1888)* 3091(1870)* ; 3093(2156)
g1957 or 4197(1921)* 4196(1605)* ; 4198(2157)
g1958 or 3121(1894)* 3120(1871)* ; 3122(2158)
g1959 or 4179(1608)* 4178(1872)* ; 4180(2159)
g1960 or 3526(1610)* 3525(1873)* ; 3527(2160)
g1961 and 845(980) 805(1844) ; 941(2161)
g1962 and 845(980) 805(1844) ; 937(2162)
g1963 and 845(980) 792(1841) 805(1844) ; 926(2163)
g1964 and 1068(981) 1038(1843) ; 1132(2164)
g1965 and 1068(981) 1026(1842) 1038(1843) ; 1126(2165)
g1966 and 827(1874) ; 5162(2166)
g1967 and 827(1874) ; 5074(2167)
g1968 and 1055(1875) ; 4780(2168)
g1969 and 3200(982) 3176(1840) 3186(1845) ; 3232(2169)
g1970 or 4316(1899)* 4315(1877)* ; 4317(2170)
g1971 or 4220(1619)* 4219(1942)* ; 4221(2171)
g1972 or 3567(1878)* 3566(1940)* ; 3568(2172)
g1973 or 4290(1911)* 4289(1880)* ; 4291(2173)
g1974 or 3535(1885)* 3534(1882)* ; 3536(2174)
g1975 or 3109(1892)* 3108(1883)* ; 3110(2175)
g1976 or 4188(1887)* 4187(1884)* ; 4189(2176)
g1977 or 3101(1907)* 3100(1886)* ; 3102(2177)
g1978 or 4594(1890)* 4593(1889)* ; 4595(2178)
g1979 or 3081(1641)* 3080(1920)* ; 3082(2179)
g1980 or 3118(1644)* 3117(1930)* ; 3119(2180)
g1981 or 7584(1906)* 7583(1891)* ; 7614(2181)
g1982 or 4585(1908)* 4584(1893)* ; 4586(2182)
g1983 or 4576(1650)* 4575(1909)* ; 4577(2183)
g1984 or 4562(1895)* 4561(1897)* ; 4563(2184)
g1985 or 4335(1653)* 4334(1939)* ; 4336(2185)
g1986 or 4326(1655)* 4325(1941)* ; 4327(2186)
g1987 or 4571(1898)* 4570(1896)* ; 4572(2187)
g1988 or 4343(1658)* 4342(1936)* ; 4344(2188)
g1989 not 4554(1900) ; 4558(2189)
g1990 or 6764(1901)* 6763(1918)* ; 6809(2190)
g1991 not 7337(1902) ; 7343(2191)
g1992 or 3051(1669)* 3050(1903)* ; 3052(2192)
g1993 or 7594(1904)* 7593(1905)* ; 7611(2193)
g1994 or 3061(1672)* 3060(1919)* ; 3062(2194)
g1995 or 3070(1675)* 3069(1934)* ; 3071(2195)
g1996 or 7550(1910)* 7549(1913)* ; 7603(2196)
g1997 or 7540(1914)* 7539(1916)* ; 7606(2197)
g1998 not 4203(1923) ; 4207(2198)
g1999 or 3549(1696)* 3548(1924)* ; 3550(2199)
g2000 or 4977(1835)* 4970(718)* ; 4979(2200)
g2001 not 1154(1928) ; 1155(2201)
g2002 or 4936(1834)* 4929(564)* ; 4938(2202)
g2003 not 7340(1931) ; 7344(2203)
g2004 or 6754(1933)* 6753(1932)* ; 6812(2204)
g2005 or 3558(1938)* 3557(1935)* ; 3559(2205)
g2006 not 4212(1937) ; 4216(2206)
g2007 or 4354(1943)* 4353(1720)* ; 4355(2207)
g2008 not 6261(1944) ; 6267(2208)
g2009 or 5936(1949)* 5929(1048)* ; 2471(2209)
g2010 or 6056(1948)* 6049(1049)* ; 2741(2210)
g2011 not 1240(1950) ; 1244(2211)
g2012 and 1258(1951) ; 1296(2212)
g2013 and 1258(1951) ; 1292(2213)
g2014 not 1249(1952) ; 1253(2214)
g2015 not 7353(1954) ; 7359(2215)
g2016 not 7356(1955) ; 7360(2216)
g2017 not 5362(1956) ; 5366(2217)
g2018 not 5359(1957) ; 5365(2218)
g2019 and 1235(1958) ; 1288(2219)
g2020 and 1235(1958) ; 1284(2220)
g2021 not 1226(1959) ; 1230(2221)
g2022 not 1217(1960) ; 1221(2222)
g2023 and 3228(2097) 3216(1462) ; 3249(2223)
g2024 and 3845(1963) 3856(1966) 3874(1968) 3989(1969) ; 4004(2224)
g2025 and 3845(1963) ; 7026(2225)
g2026 and 3845(1963) ; 6968(2226)
g2027 and 3283(1964) ; 6642(2227)
g2028 and 3283(1964) ; 6650(2228)
g2029 and 3283(1964) 3314(1967) 3344(1970) 3295(1965) ; 3431(2229)
g2030 and 3308(1109) 3283(1964) ; 3434(2230)
g2031 and 3868(1110) 3845(1963) ; 4007(2231)
g2032 and 3295(1965) ; 6666(2232)
g2033 and 3295(1965) ; 6658(2233)
g2034 and 3295(1965) 3314(1967) 3344(1970) ; 3440(2234)
g2035 and 3856(1966) ; 6978(2235)
g2036 and 3856(1966) 3874(1968) 3989(1969) ; 4013(2236)
g2037 and 3856(1966) ; 7036(2237)
g2038 and 3327(1111) 3283(1964) 3295(1965) ; 3435(2238)
g2039 and 3327(1111) 3295(1965) ; 3438(2239)
g2040 and 3327(1111) 3295(1965) ; 3441(2240)
g2041 and 3885(1112) 3856(1966) ; 4014(2241)
g2042 and 3885(1112) 3845(1963) 3856(1966) ; 4008(2242)
g2043 and 3885(1112) 3856(1966) ; 4011(2243)
g2044 and 3314(1967) ; 6682(2244)
g2045 and 3314(1967) ; 6674(2245)
g2046 and 3314(1967) 3344(1970) ; 3444(2246)
g2047 and 3874(1968) 3989(1969) ; 4051(2247)
g2048 and 3874(1968) ; 6958(2248)
g2049 and 3874(1968) ; 7016(2249)
g2050 and 3295(1965) 3335(1113) 3283(1964) 3314(1967) ; 3436(2250)
g2051 and 3295(1965) 3314(1967) 3335(1113) ; 3442(2251)
g2052 and 3295(1965) 3335(1113) 3314(1967) ; 3439(2252)
g2053 and 3335(1113) 3314(1967) ; 3443(2253)
g2054 and 3335(1113) 3314(1967) ; 3445(2254)
g2055 and 3856(1966) 3891(1114) 3874(1968) ; 4012(2255)
g2056 and 3856(1966) 3891(1114) 3845(1963) 3874(1968) ; 4009(2256)
g2057 and 3856(1966) 3891(1114) 3874(1968) ; 4015(2257)
g2058 and 3891(1114) 3874(1968) ; 4016(2258)
g2059 and 3989(1969) ; 7006(2259)
g2060 and 3989(1969) ; 6948(2260)
g2061 not 3344(1970) ; 3350(2261)
g2062 and 3899(1971) ; 7182(2262)
g2063 and 3899(1971) ; 7094(2263)
g2064 and 3899(1971) 3911(1974) 3932(1975) 3957(1977) 3997(1980) ; 4020(2264)
g2065 and 3399(1978) 3353(1972) 3381(1976) 3417(1979) 3365(1973) ; 3446(2265)
g2066 and 3353(1972) ; 4804(2266)
g2067 and 3376(1119) 3353(1972) ; 3449(2267)
g2068 and 3926(1120) 3899(1971) ; 4024(2268)
g2069 and 3365(1973) ; 4812(2269)
g2070 and 3911(1974) ; 7124(2270)
g2071 and 3957(1977) 3911(1974) 3932(1975) 3997(1980) ; 4038(2271)
g2072 and 3911(1974) ; 7114(2272)
g2073 and 3393(1121) 3365(1973) ; 3456(2273)
g2074 and 3393(1121) 3353(1972) 3365(1973) ; 3450(2274)
g2075 and 3949(1122) 3911(1974) ; 4039(2275)
g2076 and 3949(1122) 3911(1974) ; 4035(2276)
g2077 and 3949(1122) 3899(1971) 3911(1974) ; 4025(2277)
g2078 and 3932(1975) ; 7192(2278)
g2079 and 3932(1975) ; 7104(2279)
g2080 and 3957(1977) 3932(1975) 3997(1980) ; 4044(2280)
g2081 and 3381(1976) ; 4820(2281)
g2082 and 3365(1973) 3410(1123) 3381(1976) ; 3457(2282)
g2083 and 3365(1973) 3410(1123) 3353(1972) 3381(1976) ; 3451(2283)
g2084 and 3381(1976) 3410(1123) ; 3460(2284)
g2085 and 3911(1974) 3971(1124) 3932(1975) ; 4040(2285)
g2086 and 3911(1974) 3971(1124) 3932(1975) ; 4036(2286)
g2087 and 3911(1974) 3971(1124) 3899(1971) 3932(1975) ; 4026(2287)
g2088 and 3971(1124) 3932(1975) ; 4045(2288)
g2089 and 3971(1124) 3932(1975) ; 4042(2289)
g2090 and 3957(1977) ; 7084(2290)
g2091 and 3957(1977) ; 7172(2291)
g2092 and 3957(1977) 3997(1980) ; 4052(2292)
g2093 and 3399(1978) ; 4828(2293)
g2094 and 3365(1973) 3425(1125) 3381(1976) 3399(1978) ; 3458(2294)
g2095 and 3365(1973) 3425(1125) 3353(1972) 3381(1976) 3399(1978) ; 3452(2295)
g2096 and 3425(1125) 3399(1978) ; 3463(2296)
g2097 and 3425(1125) 3381(1976) 3399(1978) ; 3461(2297)
g2098 and 3911(1974) 3979(1126) 3932(1975) 3957(1977) ; 4037(2298)
g2099 and 3911(1974) 3979(1126) 3899(1971) 3932(1975) 3957(1977) ; 4027(2299)
g2100 and 3911(1974) 3979(1126) 3932(1975) 3957(1977) ; 4041(2300)
g2101 and 3979(1126) 3932(1975) 3957(1977) ; 4043(2301)
g2102 and 3979(1126) 3957(1977) ; 4047(2302)
g2103 and 3979(1126) 3932(1975) 3957(1977) ; 4046(2303)
g2104 and 3417(1979) ; 4796(2304)
g2105 and 3997(1980) ; 7162(2305)
g2106 and 3997(1980) ; 7074(2306)
g2107 and 2589(1981) 2600(1984) 2618(1985) 2734(1987) ; 2749(2307)
g2108 and 2589(1981) ; 6158(2308)
g2109 and 2589(1981) ; 6100(2309)
g2110 and 2343(1982) ; 5940(2310)
g2111 and 2343(1982) ; 5948(2311)
g2112 and 2343(1982) 2372(1986) 2400(1988) 2354(1983) ; 2487(2312)
g2113 and 2366(1130) 2343(1982) ; 2492(2313)
g2114 and 2612(1131) 2589(1981) ; 2754(2314)
g2115 and 2354(1983) ; 5964(2315)
g2116 and 2354(1983) ; 5956(2316)
g2117 and 2354(1983) 2372(1986) 2400(1988) ; 2502(2317)
g2118 and 2600(1984) ; 6110(2318)
g2119 and 2600(1984) 2618(1985) 2734(1987) ; 2764(2319)
g2120 and 2600(1984) ; 6168(2320)
g2121 and 2384(1132) 2343(1982) 2354(1983) ; 2493(2321)
g2122 and 2384(1132) 2354(1983) ; 2500(2322)
g2123 and 2384(1132) 2354(1983) ; 2503(2323)
g2124 and 2629(1133) 2600(1984) ; 2765(2324)
g2125 and 2629(1133) 2589(1981) 2600(1984) ; 2755(2325)
g2126 and 2629(1133) 2600(1984) ; 2762(2326)
g2127 and 2618(1985) 2734(1987) ; 2804(2327)
g2128 and 2618(1985) ; 6090(2328)
g2129 and 2618(1985) ; 6148(2329)
g2130 and 2372(1986) ; 5980(2330)
g2131 and 2372(1986) ; 5972(2331)
g2132 and 2372(1986) 2400(1988) ; 2506(2332)
g2133 and 2354(1983) 2391(1134) 2343(1982) 2372(1986) ; 2494(2333)
g2134 and 2354(1983) 2372(1986) 2391(1134) ; 2504(2334)
g2135 and 2354(1983) 2391(1134) 2372(1986) ; 2501(2335)
g2136 and 2391(1134) 2372(1986) ; 2505(2336)
g2137 and 2391(1134) 2372(1986) ; 2507(2337)
g2138 and 2600(1984) 2635(1135) 2618(1985) ; 2763(2338)
g2139 and 2600(1984) 2635(1135) 2589(1981) 2618(1985) ; 2756(2339)
g2140 and 2600(1984) 2635(1135) 2618(1985) ; 2766(2340)
g2141 and 2635(1135) 2618(1985) ; 2767(2341)
g2142 and 2734(1987) ; 6138(2342)
g2143 and 2734(1987) ; 6080(2343)
g2144 not 2400(1988) ; 2406(2344)
g2145 and 2409(1989) ; 4844(2345)
g2146 and 2643(1990) ; 6314(2346)
g2147 and 2643(1990) ; 6226(2347)
g2148 and 2431(1140) 2409(1989) ; 2511(2348)
g2149 and 2670(1141) 2643(1990) ; 2776(2349)
g2150 and 2655(1991) ; 6256(2350)
g2151 and 2655(1991) ; 6246(2351)
g2152 and 2420(1992) ; 4852(2352)
g2153 and 2448(1142) 2420(1992) ; 2518(2353)
g2154 and 2448(1142) 2409(1989) 2420(1992) ; 2512(2354)
g2155 and 2693(1143) 2655(1991) ; 2792(2355)
g2156 and 2693(1143) 2655(1991) ; 2788(2356)
g2157 and 2693(1143) 2643(1990) 2655(1991) ; 2777(2357)
g2158 and 2436(1993) ; 4860(2358)
g2159 and 2676(1994) ; 6324(2359)
g2160 and 2676(1994) ; 6236(2360)
g2161 and 2420(1992) 2465(1144) 2436(1993) ; 2519(2361)
g2162 and 2420(1992) 2465(1144) 2409(1989) 2436(1993) ; 2513(2362)
g2163 and 2436(1993) 2465(1144) ; 2523(2363)
g2164 and 2655(1991) 2715(1145) 2676(1994) ; 2793(2364)
g2165 and 2655(1991) 2715(1145) 2676(1994) ; 2789(2365)
g2166 and 2655(1991) 2715(1145) 2643(1990) 2676(1994) ; 2778(2366)
g2167 and 2715(1145) 2676(1994) ; 2798(2367)
g2168 and 2715(1145) 2676(1994) ; 2795(2368)
g2169 and 2701(1995) ; 6216(2369)
g2170 and 2701(1995) ; 6304(2370)
g2171 and 2454(1996) ; 4868(2371)
g2172 or 3027(2040) 3026(2020) 3025(2005) 2962(867) ; 3028(2372)
g2173 or 7602(2021)* 7595(1801)* ; 7437(2373)
g2174 and 3029(2043) 3022(1998) ; 3035(2374)
g2175 and 1718(2046) 1702(1999) ; 1788(2375)
g2176 not 5566(2000) ; 5570(2376)
g2177 not 5508(2001) ; 5512(2377)
g2178 or 1707(2029) 1706(2015) 1705(2010) 1553(870) ; 1708(2378)
g2179 or 1940(2032) 1939(2017) 1938(2006) 1802(871) ; 1941(2379)
g2180 not 5820(2002) ; 5824(2380)
g2181 not 5828(2003) ; 5832(2381)
g2182 and 1950(2047) 1935(2004) ; 1974(2382)
g2183 and 1946(2033)* 1945(2019)* 1816(875)* ; 5825(2383)
g2184 or 1944(2009) 1943(2034) 1942(2018) 1816(875) ; 5817(2384)
g2185 not 5844(2007) ; 5848(2385)
g2186 not 5836(2008) ; 5840(2386)
g2187 and 1713(2030)* 1712(2014)* 1567(876)* ; 5536(2387)
g2188 or 1711(2012) 1710(2028) 1709(2016) 1567(876) ; 5478(2388)
g2189 not 5518(2011) ; 5522(2389)
g2190 not 5576(2013) ; 5580(2390)
g2191 or 1714(2031) 1584(877) ; 1715(2391)
g2192 and 1949(2036)* 1834(878)* ; 5841(2392)
g2193 or 1948(2027) 1947(2035) 1834(878) ; 5833(2393)
g2194 or 7601(1997)* 7598(1809)* ; 7436(2394)
g2195 not 5498(2023) ; 5502(2395)
g2196 not 5556(2024) ; 5560(2396)
g2197 not 5860(2025) ; 5864(2397)
g2198 not 5852(2026) ; 5856(2398)
g2199 or 5863(1520)* 5860(2025)* ; 2003(2399)
g2200 or 5855(1161)* 5852(2026)* ; 1999(2400)
g2201 not 5546(2038) ; 5550(2401)
g2202 not 5488(2039) ; 5492(2402)
g2203 or 3033(2092) 3032(2079) 3031(2061) 3030(2055) 2989(889) ; 3034(2403)
g2204 and 4602(2041) 4535(2093) 4544(2062) ; 4626(2404)
g2205 not 4602(2041) ; 4605(2405)
g2206 not 4598(2042) ; 4601(2406)
g2207 or 1725(2081) 1724(2069) 1723(2058) 1722(2049) 1606(892) ; 1726(2407)
g2208 not 5722(2044) ; 5726(2408)
g2209 not 5634(2045) ; 5638(2409)
g2210 not 1718(2046) ; 1721(2410)
g2211 or 1956(2087) 1955(2073) 1954(2060) 1953(2050) 1866(893) ; 1957(2411)
g2212 not 4724(2048) ; 4728(2412)
g2213 and 1739(2082)* 1738(2067)* 1737(2056)* 1624(894)* ; 5692(2413)
g2214 or 1736(2053) 1735(2080) 1734(2068) 1733(2057) 1624(894) ; 5604(2414)
g2215 not 4732(2051) ; 4736(2415)
g2216 not 5664(2052) ; 5668(2416)
g2217 not 5654(2054) ; 5658(2417)
g2218 and 1744(2085)* 1743(2070)* 1647(899)* ; 5672(2418)
g2219 or 1742(2065) 1741(2083) 1740(2071) 1647(899) ; 5584(2419)
g2220 and 4598(2042) 4531(1830) 4540(1822) ; 4623(2420)
g2221 not 5732(2063) ; 5736(2421)
g2222 not 5644(2064) ; 5648(2422)
g2223 not 4740(2066) ; 4744(2423)
g2224 or 1745(2084) 1669(904) ; 1746(2424)
g2225 not 4748(2075) ; 4752(2425)
g2226 not 5624(2076) ; 5628(2426)
g2227 not 5712(2077) ; 5716(2427)
g2228 not 5702(2090) ; 5706(2428)
g2229 not 5614(2091) ; 5618(2429)
g2230 not 4716(2094) ; 4720(2430)
g2231 and 1122(2101) 1108(1196) ; 1146(2431)
g2232 and 920(2100) 902(1199) ; 997(2432)
g2233 or 928(2126) 927(2112) 926(2163) 925(2103) 802(924) ; 929(2433)
g2234 or 1128(2132) 1127(2116) 1126(2165) 1125(2104) 1035(925) ; 1129(2434)
g2235 or 3234(2137) 3233(2119) 3232(2169) 3231(2109) 3183(926) ; 3235(2435)
g2236 and 3575(2095) 3508(2138) 3517(2120) ; 3599(2436)
g2237 not 3575(2095) ; 3578(2437)
g2238 not 3571(2096) ; 3574(2438)
g2239 not 5152(2098) ; 5156(2439)
g2240 not 5064(2099) ; 5068(2440)
g2241 not 920(2100) ; 924(2441)
g2242 not 4764(2102) ; 4768(2442)
g2243 and 943(2127)* 942(2110)* 941(2161)* 821(929)* ; 5122(2443)
g2244 or 940(2107) 939(2125) 938(2111) 937(2162) 821(929) ; 5034(2444)
g2245 not 4772(2105) ; 4776(2445)
g2246 not 5094(2106) ; 5098(2446)
g2247 not 5084(2108) ; 5088(2447)
g2248 or 949(2129) 868(934) ; 950(2448)
g2249 not 4788(2118) ; 4792(2449)
g2250 and 3571(2096) 3504(1851) 3513(1848) ; 3596(2450)
g2251 not 5054(2121) ; 5058(2451)
g2252 not 5142(2123) ; 5146(2452)
g2253 not 5132(2135) ; 5136(2453)
g2254 not 5044(2136) ; 5048(2454)
g2255 not 4756(2139) ; 4760(2455)
g2256 and 4263(2142) 4226(1854) 4235(1855) ; 4284(2456)
g2257 and 4267(2143) 4230(2140) 4239(2141) ; 4287(2457)
g2258 not 4263(2142) ; 4266(2458)
g2259 not 4267(2143) ; 4270(2459)
g2260 and 1300(2146) 1263(1857) 1272(1858) ; 1321(2460)
g2261 and 1304(2147) 1267(2144) 1276(2145) ; 1324(2461)
g2262 not 1300(2146) ; 1303(2462)
g2263 not 1304(2147) ; 1307(2463)
g2264 not 7348(2148) ; 7352(2464)
g2265 and 4300(2153) 4314(1248) 4291(2173) 4308(2151) ; 4363(2465)
g2266 and 4291(2173) 4300(2153) 4308(2151) 4352(2149) ; 4356(2466)
g2267 not 6822(2150) ; 6826(2467)
g2268 and 4312(1256) 4291(2173) 4300(2153) ; 4362(2468)
g2269 not 6819(2152) ; 6825(2469)
g2270 and 4305(1262) 4291(2173) ; 4361(2470)
g2271 not 7345(2154) ; 7351(2471)
g2272 and 3545(2155) ; 3583(2472)
g2273 and 3545(2155) ; 3579(2473)
g2274 and 3099(1268) 3082(2179) ; 3139(2474)
g2275 and 3082(2179) 3093(2156) 3102(2177) 3110(2175) 3122(2158) ; 3136(2475)
g2276 and 4198(2157) ; 4251(2476)
g2277 and 4198(2157) ; 4247(2477)
g2278 and 3093(2156) 3116(1271) 3082(2179) 3102(2177) 3110(2175) ; 3142(2478)
g2279 not 4180(2159) ; 4184(2479)
g2280 not 3527(2160) ; 3531(2480)
g2281 and 948(2130)* 947(2113)* 845(980)* ; 5102(2481)
g2282 or 946(2122) 945(2128) 944(2114) 845(980) ; 5014(2482)
g2283 not 5162(2166) ; 5166(2483)
g2284 not 5074(2167) ; 5078(2484)
g2285 not 4780(2168) ; 4784(2485)
g2286 and 4317(2170) 4327(2186) 4336(2185) 4344(2188) 4355(2207) ; 4369(2486)
g2287 and 4221(2171) ; 4259(2487)
g2288 and 4221(2171) ; 4255(2488)
g2289 and 3568(2172) ; 3587(2489)
g2290 and 3568(2172) ; 3591(2490)
g2291 not 3536(2174) ; 3540(2491)
g2292 and 3093(2156) 3114(1298) 3082(2179) 3102(2177) ; 3141(2492)
g2293 not 4189(2176) ; 4193(2493)
g2294 and 3107(1305) 3082(2179) 3093(2156) ; 3140(2494)
g2295 and 4595(2178) ; 4614(2495)
g2296 and 4595(2178) ; 4618(2496)
g2297 and 3052(2192) 3062(2194) 3071(2195) 3119(2180) ; 3123(2497)
g2298 not 7614(2181) ; 7618(2498)
g2299 not 4586(2182) ; 4590(2499)
g2300 not 4577(2183) ; 4581(2500)
g2301 not 4563(2184) ; 4567(2501)
g2302 and 4572(2187) ; 4610(2502)
g2303 and 4572(2187) ; 4606(2503)
g2304 not 6809(2190) ; 6815(2504)
g2305 or 7344(2203)* 7337(1902)* ; 6351(2505)
g2306 not 7611(2193) ; 7617(2506)
g2307 not 7603(2196) ; 7609(2507)
g2308 not 7606(2197) ; 7610(2508)
g2309 and 3068(1353) 3052(2192) ; 3128(2509)
g2310 not 3550(2199) ; 3554(2510)
g2311 or 4979(2200)* 4978(1926)* ; 4980(2511)
g2312 or 4938(2202)* 4937(1929)* ; 4939(2512)
g2313 and 3062(2194) 3079(1370) 3052(2192) 3071(2195) ; 3130(2513)
g2314 or 7343(2191)* 7340(1931)* ; 6350(2514)
g2315 not 6812(2204) ; 6816(2515)
g2316 and 3076(1379) 3052(2192) 3062(2194) ; 3129(2516)
g2317 not 3559(2205) ; 3563(2517)
g2318 and 4327(2186) 4348(1385) 4317(2170) 4336(2185) ; 4374(2518)
g2319 and 4341(1392) 4317(2170) 4327(2186) ; 4373(2519)
g2320 and 4333(1397) 4317(2170) ; 4372(2520)
g2321 and 4327(2186) 4349(1400) 4317(2170) 4336(2185) 4344(2188) ; 4375(2521)
g2322 and 2420(1992) 2481(1721) 2436(1993) 2454(1996) ; 2520(2522)
g2323 and 2420(1992) 2481(1721) 2409(1989) 2436(1993) 2454(1996) ; 2514(2523)
g2324 and 2481(1721) 2454(1996) ; 2527(2524)
g2325 and 2481(1721) 2436(1993) 2454(1996) ; 2524(2525)
g2326 and 2655(1991) 2724(1722) 2676(1994) 2701(1995) ; 2790(2526)
g2327 and 2655(1991) 2724(1722) 2643(1990) 2676(1994) 2701(1995) ; 2779(2527)
g2328 and 2655(1991) 2724(1722) 2676(1994) 2701(1995) ; 2794(2528)
g2329 and 2724(1722) 2676(1994) 2701(1995) ; 2796(2529)
g2330 and 2724(1722) 2701(1995) ; 2800(2530)
g2331 and 2724(1722) 2676(1994) 2701(1995) ; 2799(2531)
g2332 or 2471(2209)* 2470(1945)* ; 2472(2532)
g2333 or 2741(2210)* 2740(1947)* ; 2742(2533)
g2334 and 1292(2213) 1240(1950) 1249(1952) ; 1315(2534)
g2335 and 1296(2212) 1244(2211) 1253(2214) ; 1318(2535)
g2336 not 1296(2212) ; 1299(2536)
g2337 not 1292(2213) ; 1295(2537)
g2338 or 7360(2216)* 7353(1954)* ; 6341(2538)
g2339 or 7359(2215)* 7356(1955)* ; 6340(2539)
g2340 or 5365(2218)* 5362(1956)* ; 5367(2540)
g2341 or 5366(2217)* 5359(1957)* ; 5368(2541)
g2342 and 1288(2219) 1221(2222) 1230(2221) ; 1312(2542)
g2343 not 1288(2219) ; 1291(2543)
g2344 not 1284(2220) ; 1287(2544)
g2345 and 1284(2220) 1217(1960) 1226(1959) ; 1309(2545)
g2346 and 3235(2435) 3216(1462) ; 3258(2546)
g2347 and 2472(2532) 4526(205) ; 2531(2547)
g2348 and 2454(1996) 2472(2532) 4526(205) ; 2529(2548)
g2349 and 2454(1996) 2436(1993) 2472(2532) 4526(205) ; 2526(2549)
g2350 and 2420(1992) 2454(1996) 2436(1993) 2472(2532) 4526(205) ; 2522(2550)
g2351 or 3436(2250) 3435(2238) 3434(2230) 3292(1107) ; 3437(2551)
g2352 or 4009(2256) 4008(2242) 4007(2231) 3853(1108) ; 4010(2552)
g2353 and 4020(2264) 4004(2224) ; 4089(2553)
g2354 not 7026(2225) ; 7030(2554)
g2355 not 6968(2226) ; 6972(2555)
g2356 not 6642(2227) ; 6646(2556)
g2357 not 6650(2228) ; 6654(2557)
g2358 and 3446(2265) 3431(2229) ; 3466(2558)
g2359 and 3442(2251)* 3441(2240)* 3308(1109)* ; 6647(2559)
g2360 or 3440(2234) 3439(2252) 3438(2239) 3308(1109) ; 6639(2560)
g2361 and 4015(2257)* 4014(2241)* 3868(1110)* ; 6996(2561)
g2362 or 4013(2236) 4012(2255) 4011(2243) 3868(1110) ; 6938(2562)
g2363 not 6666(2232) ; 6670(2563)
g2364 not 6658(2233) ; 6662(2564)
g2365 not 6978(2235) ; 6982(2565)
g2366 not 7036(2237) ; 7040(2566)
g2367 and 3445(2254)* 3327(1111)* ; 6663(2567)
g2368 or 3444(2246) 3443(2253) 3327(1111) ; 6655(2568)
g2369 or 4016(2258) 3885(1112) ; 4017(2569)
g2370 not 6682(2244) ; 6686(2570)
g2371 not 6674(2245) ; 6678(2571)
g2372 not 6958(2248) ; 6962(2572)
g2373 not 7016(2249) ; 7020(2573)
g2374 or 6685(1768)* 6682(2244)* ; 3487(2574)
g2375 not 7006(2259) ; 7010(2575)
g2376 not 6948(2260) ; 6952(2576)
g2377 or 6677(1474)* 6674(2245)* ; 3483(2577)
g2378 or 3452(2295) 3451(2283) 3450(2274) 3449(2267) 3362(1117) ; 3453(2578)
g2379 or 4027(2299) 4026(2287) 4025(2277) 4024(2268) 3908(1118) ; 4028(2579)
g2380 not 7182(2262) ; 7186(2580)
g2381 not 7094(2263) ; 7098(2581)
g2382 not 4020(2264) ; 4023(2582)
g2383 not 4804(2266) ; 4808(2583)
g2384 and 4041(2300)* 4040(2285)* 4039(2275)* 3926(1120)* ; 7152(2584)
g2385 or 4038(2271) 4037(2298) 4036(2286) 4035(2276) 3926(1120) ; 7064(2585)
g2386 not 4812(2269) ; 4816(2586)
g2387 not 7124(2270) ; 7128(2587)
g2388 not 7114(2272) ; 7118(2588)
g2389 and 4046(2303)* 4045(2288)* 3949(1122)* ; 7132(2589)
g2390 or 4044(2280) 4043(2301) 4042(2289) 3949(1122) ; 7044(2590)
g2391 not 7192(2278) ; 7196(2591)
g2392 not 7104(2279) ; 7108(2592)
g2393 not 4820(2281) ; 4824(2593)
g2394 or 4047(2302) 3971(1124) ; 4048(2594)
g2395 not 7084(2290) ; 7088(2595)
g2396 not 7172(2291) ; 7176(2596)
g2397 not 4828(2293) ; 4832(2597)
g2398 not 4796(2304) ; 4800(2598)
g2399 not 7162(2305) ; 7166(2599)
g2400 not 7074(2306) ; 7078(2600)
g2401 or 2494(2333) 2493(2321) 2492(2313) 2351(1128) ; 2495(2601)
g2402 or 2756(2339) 2755(2325) 2754(2314) 2597(1129) ; 2757(2602)
g2403 not 2749(2307) ; 2753(2603)
g2404 not 6158(2308) ; 6162(2604)
g2405 not 6100(2309) ; 6104(2605)
g2406 not 5940(2310) ; 5944(2606)
g2407 not 5948(2311) ; 5952(2607)
g2408 not 2487(2312) ; 2491(2608)
g2409 and 2504(2334)* 2503(2323)* 2366(1130)* ; 5945(2609)
g2410 or 2502(2317) 2501(2335) 2500(2322) 2366(1130) ; 5937(2610)
g2411 and 2766(2340)* 2765(2324)* 2612(1131)* ; 6128(2611)
g2412 or 2764(2319) 2763(2338) 2762(2326) 2612(1131) ; 6070(2612)
g2413 not 5964(2315) ; 5968(2613)
g2414 not 5956(2316) ; 5960(2614)
g2415 not 6110(2318) ; 6114(2615)
g2416 not 6168(2320) ; 6172(2616)
g2417 and 2507(2337)* 2384(1132)* ; 5961(2617)
g2418 or 2506(2332) 2505(2336) 2384(1132) ; 5953(2618)
g2419 or 2767(2341) 2629(1133) ; 2768(2619)
g2420 not 6090(2328) ; 6094(2620)
g2421 not 6148(2329) ; 6152(2621)
g2422 not 5980(2330) ; 5984(2622)
g2423 not 5972(2331) ; 5976(2623)
g2424 or 5983(1789)* 5980(2330)* ; 2559(2624)
g2425 not 6138(2342) ; 6142(2625)
g2426 not 6080(2343) ; 6084(2626)
g2427 or 5975(1498)* 5972(2331)* ; 2555(2627)
g2428 or 2514(2523) 2513(2362) 2512(2354) 2511(2348) 2417(1138) ; 2515(2628)
g2429 or 2779(2527) 2778(2366) 2777(2357) 2776(2349) 2652(1139) ; 2780(2629)
g2430 and 2454(1996) 2409(1989) 2436(1993) 2472(2532) 2420(1992) ; 2508(2630)
g2431 not 4844(2345) ; 4848(2631)
g2432 not 6314(2346) ; 6318(2632)
g2433 not 6226(2347) ; 6230(2633)
g2434 and 2643(1990) 2655(1991) 2676(1994) 2701(1995) 2742(2533) ; 2771(2634)
g2435 and 2794(2528)* 2793(2364)* 2792(2355)* 2670(1141)* ; 6284(2635)
g2436 not 6256(2350) ; 6260(2636)
g2437 and 2701(1995) 2655(1991) 2676(1994) 2742(2533) ; 2791(2637)
g2438 not 6246(2351) ; 6250(2638)
g2439 not 4852(2352) ; 4856(2639)
g2440 and 2799(2531)* 2798(2367)* 2693(1143)* ; 6264(2640)
g2441 not 4860(2358) ; 4864(2641)
g2442 not 6324(2359) ; 6328(2642)
g2443 not 6236(2360) ; 6240(2643)
g2444 and 2701(1995) 2676(1994) 2742(2533) ; 2797(2644)
g2445 or 2800(2530) 2715(1145) ; 2801(2645)
g2446 not 6216(2369) ; 6220(2646)
g2447 not 6304(2370) ; 6308(2647)
g2448 and 2701(1995) 2742(2533) ; 2807(2648)
g2449 not 4868(2371) ; 4872(2649)
g2450 or 7437(2373)* 7436(2394)* ; 7438(2650)
g2451 and 3034(2403) 3022(1998) ; 3045(2651)
g2452 and 1726(2407) 1702(1999) ; 1789(2652)
g2453 or 5824(2380)* 5817(2384)* ; 1986(2653)
g2454 or 5832(2381)* 5825(2383)* ; 1989(2654)
g2455 and 1935(2004) 1957(2411) ; 1981(2655)
g2456 not 5825(2383) ; 5831(2656)
g2457 not 5817(2384) ; 5823(2657)
g2458 or 5848(2385)* 5841(2392)* ; 1996(2658)
g2459 or 5840(2386)* 5833(2393)* ; 1993(2659)
g2460 not 5536(2387) ; 5540(2660)
g2461 not 5478(2388) ; 5482(2661)
g2462 not 1715(2391) ; 5526(2662)
g2463 not 5841(2392) ; 5847(2663)
g2464 not 5833(2393) ; 5839(2664)
g2465 or 1749(2022) 1715(2391) ; 5468(2665)
g2466 or 5864(2397)* 5857(1159)* ; 2004(2666)
g2467 or 5856(2398)* 5849(884)* ; 2000(2667)
g2468 not 1726(2407) ; 1730(2668)
g2469 not 5692(2413) ; 5696(2669)
g2470 not 5604(2414) ; 5608(2670)
g2471 not 5672(2418) ; 5676(2671)
g2472 not 5584(2419) ; 5588(2672)
g2473 and 4601(2406) 4540(1822) 4535(2093) ; 4622(2673)
g2474 not 1746(2424) ; 5682(2674)
g2475 or 1750(2078) 1746(2424) ; 5594(2675)
g2476 or 5675(1541)* 5672(2418)* ; 5677(2676)
g2477 or 5587(1183)* 5584(2419)* ; 5589(2677)
g2478 and 4605(2405) 4544(2062) 4531(1830) ; 4625(2678)
g2479 or 4987(1549)* 4980(2511)* ; 4989(2679)
g2480 or 4946(1837)* 4939(2512)* ; 4948(2680)
g2481 and 1108(1196) 1129(2434) ; 1151(2681)
g2482 and 929(2433) 902(1199) ; 1002(2682)
g2483 not 929(2433) ; 933(2683)
g2484 not 3235(2435) ; 3238(2684)
g2485 not 5122(2443) ; 5126(2685)
g2486 not 5034(2444) ; 5038(2686)
g2487 not 950(2448) ; 5112(2687)
g2488 and 3574(2438) 3513(1848) 3508(2138) ; 3595(2688)
g2489 or 956(2124) 950(2448) ; 5024(2689)
g2490 or 5105(1569)* 5102(2481)* ; 5107(2690)
g2491 or 5017(1219)* 5014(2482)* ; 5019(2691)
g2492 and 3578(2437) 3517(2120) 3504(1851) ; 3598(2692)
g2493 and 4270(2459) 4239(2141) 4226(1854) ; 4286(2693)
g2494 and 4266(2458) 4235(1855) 4230(2140) ; 4283(2694)
g2495 and 1307(2463) 1276(2145) 1263(1857) ; 1323(2695)
g2496 and 1303(2462) 1272(1858) 1267(2144) ; 1320(2696)
g2497 or 7351(2471)* 7348(2148)* ; 6360(2697)
g2498 and 4369(2486) 4356(2466) ; 4386(2698)
g2499 not 4356(2466) ; 4360(2699)
g2500 or 6825(2469)* 6822(2150)* ; 6827(2700)
g2501 or 6826(2467)* 6819(2152)* ; 6828(2701)
g2502 or 7352(2464)* 7345(2154)* ; 6361(2702)
g2503 and 3583(2472) 3531(2480) 3540(2491) ; 3605(2703)
g2504 not 3583(2472) ; 3586(2704)
g2505 not 3579(2473) ; 3582(2705)
g2506 and 3136(2475) 3123(2497) ; 3156(2706)
g2507 and 4251(2476) 4184(2479) 4193(2493) ; 4275(2707)
g2508 not 4251(2476) ; 4254(2708)
g2509 not 4247(2477) ; 4250(2709)
g2510 and 4247(2477) 4180(2159) 4189(2176) ; 4272(2710)
g2511 and 3579(2473) 3527(2160) 3536(2174) ; 3602(2711)
g2512 not 5102(2481) ; 5106(2712)
g2513 not 5014(2482) ; 5018(2713)
g2514 or 4375(2521) 4374(2518) 4373(2519) 4372(2520) 4324(1284) ; 4376(2714)
g2515 not 4259(2487) ; 4262(2715)
g2516 not 4255(2488) ; 4258(2716)
g2517 not 3587(2489) ; 3590(2717)
g2518 and 3591(2490) 3554(2510) 3563(2517) ; 3611(2718)
g2519 not 3591(2490) ; 3594(2719)
g2520 or 4363(2465) 4362(2468) 4361(2470) 4297(1293) ; 4364(2720)
g2521 or 89(48)* 4369(2486)* ; 4380(2721)
g2522 not 4614(2495) ; 4617(2722)
g2523 and 4618(2496) 4581(2500) 4590(2499) ; 4638(2723)
g2524 not 4618(2496) ; 4621(2724)
g2525 not 3123(2497) ; 3127(2725)
g2526 or 7617(2506)* 7614(2181)* ; 7446(2726)
g2527 and 4614(2495) 4577(2183) 4586(2182) ; 4635(2727)
g2528 not 4610(2502) ; 4613(2728)
g2529 not 4606(2503) ; 4609(2729)
g2530 and 4606(2503) 4554(1900) 4563(2184) ; 4629(2730)
g2531 and 4610(2502) 4558(2189) 4567(2501) ; 4632(2731)
g2532 or 6816(2515)* 6809(2190)* ; 6818(2732)
g2533 or 3130(2513) 3129(2516) 3128(2509) 3059(1330) ; 3131(2733)
g2534 or 6351(2505)* 6350(2514)* ; 6352(2734)
g2535 or 7618(2498)* 7611(2193)* ; 7447(2735)
g2536 or 7610(2508)* 7603(2196)* ; 7457(2736)
g2537 or 7609(2507)* 7606(2197)* ; 7456(2737)
g2538 or 3142(2478) 3141(2492) 3140(2494) 3139(2474) 3090(1356) ; 3143(2738)
g2539 and 4255(2488) 4203(1923) 4212(1937) ; 4278(2739)
g2540 and 4259(2487) 4207(2198) 4216(2206) ; 4281(2740)
g2541 and 3587(2489) 3550(2199) 3559(2205) ; 3608(2741)
g2542 not 4980(2511) ; 4986(2742)
g2543 not 4939(2512) ; 4945(2743)
g2544 or 6815(2504)* 6812(2204)* ; 6817(2744)
g2545 and 2472(2532) ; 4836(2745)
g2546 and 2742(2533) ; 6294(2746)
g2547 and 2742(2533) ; 6206(2747)
g2548 and 1299(2536) 1253(2214) 1240(1950) ; 1317(2748)
g2549 and 1295(2537) 1249(1952) 1244(2211) ; 1314(2749)
g2550 or 6341(2538)* 6340(2539)* ; 6342(2750)
g2551 or 5368(2541)* 5367(2540)* ; 5388(2751)
g2552 and 1287(2544) 1226(1959) 1221(2222) ; 1308(2752)
g2553 and 1291(2543) 1230(2221) 1217(1960) ; 1311(2753)
g2554 or 4839(316)* 4836(2745)* ; 371(2754)
g2555 or 4526(205)* 2771(2634)* ; 2806(2755)
g2556 and 4526(205) 2508(2630) ; 2563(2756)
g2557 and 4028(2579) 4004(2224) ; 4090(2757)
g2558 or 6646(2556)* 6639(2560)* ; 3470(2758)
g2559 or 6654(2557)* 6647(2559)* ; 3473(2759)
g2560 and 3431(2229) 3453(2578) ; 3467(2760)
g2561 not 6647(2559) ; 6653(2761)
g2562 not 6639(2560) ; 6645(2762)
g2563 not 6996(2561) ; 7000(2763)
g2564 not 6938(2562) ; 6942(2764)
g2565 or 6670(2563)* 6663(2567)* ; 3480(2765)
g2566 or 6662(2564)* 6655(2568)* ; 3477(2766)
g2567 not 6663(2567) ; 6669(2767)
g2568 not 6655(2568) ; 6661(2768)
g2569 not 4017(2569) ; 6986(2769)
g2570 or 4051(2247) 4017(2569) ; 6928(2770)
g2571 or 6686(2570)* 6679(1469)* ; 3488(2771)
g2572 or 6678(2571)* 6671(1116)* ; 3484(2772)
g2573 not 4028(2579) ; 4032(2773)
g2574 not 7152(2584) ; 7156(2774)
g2575 not 7064(2585) ; 7068(2775)
g2576 not 7132(2589) ; 7136(2776)
g2577 not 7044(2590) ; 7048(2777)
g2578 not 4048(2594) ; 7142(2778)
g2579 or 4052(2292) 4048(2594) ; 7054(2779)
g2580 or 7135(1780)* 7132(2589)* ; 7137(2780)
g2581 or 7047(1485)* 7044(2590)* ; 7049(2781)
g2582 not 2495(2601) ; 2499(2782)
g2583 not 2757(2602) ; 2761(2783)
g2584 and 2780(2629) 2749(2307) ; 2853(2784)
g2585 and 2771(2634) 2749(2307) ; 2852(2785)
g2586 or 5944(2606)* 5937(2610)* ; 2542(2786)
g2587 or 5952(2607)* 5945(2609)* ; 2545(2787)
g2588 and 2508(2630) 2487(2312) ; 2532(2788)
g2589 and 2487(2312) 2515(2628) ; 2536(2789)
g2590 not 5945(2609) ; 5951(2790)
g2591 not 5937(2610) ; 5943(2791)
g2592 not 6128(2611) ; 6132(2792)
g2593 not 6070(2612) ; 6074(2793)
g2594 or 5968(2613)* 5961(2617)* ; 2552(2794)
g2595 or 5960(2614)* 5953(2618)* ; 2549(2795)
g2596 not 5961(2617) ; 5967(2796)
g2597 not 5953(2618) ; 5959(2797)
g2598 not 2768(2619) ; 6118(2798)
g2599 or 2804(2327) 2768(2619) ; 6060(2799)
g2600 or 5984(2622)* 5977(1493)* ; 2560(2800)
g2601 or 5976(2623)* 5969(1137)* ; 2556(2801)
g2602 not 2780(2629) ; 2784(2802)
g2603 not 2771(2634) ; 2775(2803)
g2604 or 2522(2550) 2520(2522) 2519(2361) 2518(2353) 2431(1140) ; 4841(2804)
g2605 not 6284(2635) ; 6288(2805)
g2606 or 2791(2637) 2790(2526) 2789(2365) 2788(2356) 2670(1141) ; 6196(2806)
g2607 or 2526(2549) 2524(2525) 2523(2363) 2448(1142) ; 4849(2807)
g2608 not 6264(2640) ; 6268(2808)
g2609 or 2797(2644) 2796(2529) 2795(2368) 2693(1143) ; 6176(2809)
g2610 or 2529(2548) 2527(2524) 2465(1144) ; 4857(2810)
g2611 or 2807(2648) 2801(2645) ; 6186(2811)
g2612 not 2801(2645) ; 6274(2812)
g2613 or 3045(2651) 3028(2372) ; 3046(2813)
g2614 not 7438(2650) ; 7442(2814)
g2615 or 1789(2652) 1708(2378) ; 1790(2815)
g2616 or 1981(2655) 1941(2379) ; 1982(2816)
g2617 or 5823(2657)* 5820(2002)* ; 1985(2817)
g2618 or 5831(2656)* 5828(2003)* ; 1988(2818)
g2619 or 5847(2663)* 5844(2007)* ; 1995(2819)
g2620 or 5839(2664)* 5836(2008)* ; 1992(2820)
g2621 not 5526(2662) ; 5530(2821)
g2622 not 5468(2665) ; 5472(2822)
g2623 or 5529(1519)* 5526(2662)* ; 5531(2823)
g2624 or 2004(2666)* 2003(2399)* ; 2005(2824)
g2625 or 2000(2667)* 1999(2400)* ; 2001(2825)
g2626 or 5471(1162)* 5468(2665)* ; 5473(2826)
g2627 and 4626(2404)* 4625(2678)* ; 4627(2827)
g2628 and 1721(2410) 1730(2668) ; 1751(2828)
g2629 and 4623(2420)* 4622(2673)* ; 4624(2829)
g2630 not 5682(2674) ; 5686(2830)
g2631 not 5594(2675) ; 5598(2831)
g2632 or 5676(2671)* 5669(1182)* ; 5678(2832)
g2633 or 5588(2672)* 5581(911)* ; 5590(2833)
g2634 or 4986(2742)* 4983(1191)* ; 4988(2834)
g2635 or 1002(2682) 908(1192) ; 265(2835)
g2636 or 4945(2743)* 4942(1551)* ; 4947(2836)
g2637 or 1151(2681) 1117(1193) ; 241(2837)
g2638 and 3599(2436)* 3598(2692)* ; 3600(2838)
g2639 and 924(2441) 933(2683) ; 962(2839)
g2640 not 5112(2687) ; 5116(2840)
g2641 and 3596(2450)* 3595(2688)* ; 3597(2841)
g2642 not 5024(2689) ; 5028(2842)
g2643 or 5106(2712)* 5099(1218)* ; 5108(2843)
g2644 or 5018(2713)* 5011(941)* ; 5020(2844)
g2645 and 4284(2456)* 4283(2694)* ; 4285(2845)
g2646 and 4287(2457)* 4286(2693)* ; 4288(2846)
g2647 and 1321(2460)* 1320(2696)* ; 1322(2847)
g2648 and 1324(2461)* 1323(2695)* ; 1325(2848)
g2649 or 6361(2702)* 6360(2697)* ; 6362(2849)
g2650 and 4376(2714) 4356(2466) ; 4387(2850)
g2651 or 6828(2701)* 6827(2700)* ; 6848(2851)
g2652 and 4254(2708) 4193(2493) 4180(2159) ; 4274(2852)
g2653 and 3586(2704) 3540(2491) 3527(2160) ; 3604(2853)
g2654 not 4376(2714) ; 4379(2854)
g2655 not 4364(2720) ; 4368(2855)
g2656 and 3582(2705) 3536(2174) 3531(2480) ; 3601(2856)
g2657 and 4250(2709) 4189(2176) 4184(2479) ; 4271(2857)
g2658 and 3249(2223) 3035(2374) 3156(2706) 4386(2698) 89(48) ; 263(2858)
g2659 and 3035(2374) 3156(2706) 4386(2698) 89(48) ; 3241(2859)
g2660 and 3249(2223) 3035(2374) 3156(2706) 4386(2698) 89(48) ; 257(2860)
g2661 and 3143(2738) 3123(2497) ; 3163(2861)
g2662 or 7447(2735)* 7446(2726)* ; 7448(2862)
g2663 and 4617(2722) 4586(2182) 4581(2500) ; 4634(2863)
g2664 and 4621(2724) 4590(2499) 4577(2183) ; 4637(2864)
g2665 and 4609(2729) 4563(2184) 4558(2189) ; 4628(2865)
g2666 and 4613(2728) 4567(2501) 4554(1900) ; 4631(2866)
g2667 or 6818(2732)* 6817(2744)* ; 6840(2867)
g2668 not 3131(2733) ; 3135(2868)
g2669 not 6352(2734) ; 6356(2869)
g2670 or 7457(2736)* 7456(2737)* ; 7458(2870)
g2671 not 3143(2738) ; 3146(2871)
g2672 and 4262(2715) 4216(2206) 4203(1923) ; 4280(2872)
g2673 and 3594(2719) 3563(2517) 3550(2199) ; 3610(2873)
g2674 or 3258(2546) 3223(1698) ; 3259(2874)
g2675 and 3590(2717) 3559(2205) 3554(2510) ; 3607(2875)
g2676 and 4258(2716) 4212(1937) 4207(2198) ; 4277(2876)
g2677 or 2531(2547) 2481(1721) ; 4865(2877)
g2678 or 6267(2208)* 6264(2640)* ; 6269(2878)
g2679 not 4836(2745) ; 4840(2879)
g2680 not 6294(2746) ; 6298(2880)
g2681 not 6206(2747) ; 6210(2881)
g2682 and 1315(2534)* 1314(2749)* ; 1316(2882)
g2683 and 1318(2535)* 1317(2748)* ; 1319(2883)
g2684 not 6342(2750) ; 6346(2884)
g2685 not 5388(2751) ; 5392(2885)
g2686 and 1312(2542)* 1311(2753)* ; 1313(2886)
g2687 and 1309(2545)* 1308(2752)* ; 1310(2887)
g2688 and 3249(2223) 3046(2813) ; 254(2888)
g2689 and 3249(2223) 3046(2813) ; 260(2889)
g2690 or 4840(2879)* 4833(207)* ; 372(2890)
g2691 and 3466(2558) 2532(2788) 4526(205) ; 3277(2891)
g2692 and 1974(2382) 3466(2558) 2532(2788) 4526(205) ; 3270(2892)
g2693 and 2806(2755) 2784(2802) ; 2809(2893)
g2694 and 4089(2553) 2852(2785) 4526(205) ; 1454(2894)
g2695 and 1788(2375) 4089(2553) 2852(2785) 4526(205) ; 1445(2895)
g2696 and 997(2432) 1788(2375) 4089(2553) 2852(2785) 4526(205) ; 269(2896)
g2697 and 1146(2431) 1974(2382) 3466(2558) 2532(2788) 4526(205) ; 245(2897)
g2698 or 3467(2760) 3437(2551) ; 3468(2898)
g2699 or 4090(2757) 4010(2552) ; 4091(2899)
g2700 or 6645(2762)* 6642(2227)* ; 3469(2900)
g2701 or 6653(2761)* 6650(2228)* ; 3472(2901)
g2702 or 6669(2767)* 6666(2232)* ; 3479(2902)
g2703 or 6661(2768)* 6658(2233)* ; 3476(2903)
g2704 not 6986(2769) ; 6990(2904)
g2705 not 6928(2770) ; 6932(2905)
g2706 or 3488(2771)* 3487(2574)* ; 3489(2906)
g2707 or 6989(1769)* 6986(2769)* ; 6991(2907)
g2708 or 6931(1471)* 6928(2770)* ; 6933(2908)
g2709 or 3484(2772)* 3483(2577)* ; 3485(2909)
g2710 and 4023(2582) 4032(2773) ; 4053(2910)
g2711 not 7142(2778) ; 7146(2911)
g2712 not 7054(2779) ; 7058(2912)
g2713 or 7136(2776)* 7129(1483)* ; 7138(2913)
g2714 or 7048(2777)* 7041(1127)* ; 7050(2914)
g2715 or 2536(2789) 2495(2601) ; 2537(2915)
g2716 or 2853(2784) 2757(2602) ; 2854(2916)
g2717 or 2753(2603)* 2761(2783)* ; 2808(2917)
g2718 or 5943(2791)* 5940(2310)* ; 2541(2918)
g2719 or 5951(2790)* 5948(2311)* ; 2544(2919)
g2720 or 2491(2608)* 2499(2782)* ; 2577(2920)
g2721 or 5967(2796)* 5964(2315)* ; 2551(2921)
g2722 or 5959(2797)* 5956(2316)* ; 2548(2922)
g2723 not 6118(2798) ; 6122(2923)
g2724 not 6060(2799) ; 6064(2924)
g2725 or 2560(2800)* 2559(2624)* ; 2561(2925)
g2726 or 6121(1790)* 6118(2798)* ; 6123(2926)
g2727 or 6063(1495)* 6060(2799)* ; 6065(2927)
g2728 or 2556(2801)* 2555(2627)* ; 2557(2928)
g2729 or 2563(2756) 2515(2628) ; 2564(2929)
g2730 and 2775(2803) 2784(2802) ; 2813(2930)
g2731 or 4848(2631)* 4841(2804)* ; 387(2931)
g2732 not 4841(2804) ; 4847(2932)
g2733 not 6196(2806) ; 6200(2933)
g2734 or 4856(2639)* 4849(2807)* ; 390(2934)
g2735 not 4849(2807) ; 4855(2935)
g2736 not 6176(2809) ; 6180(2936)
g2737 or 4864(2641)* 4857(2810)* ; 393(2937)
g2738 not 4857(2810) ; 4863(2938)
g2739 not 6186(2811) ; 6190(2939)
g2740 not 6274(2812) ; 6278(2940)
g2741 or 4872(2649)* 4865(2877)* ; 396(2941)
g2742 or 1986(2653)* 1985(2817)* ; 1987(2942)
g2743 or 1989(2654)* 1988(2818)* ; 1990(2943)
g2744 or 1996(2658)* 1995(2819)* ; 1997(2944)
g2745 or 1993(2659)* 1992(2820)* ; 1994(2945)
g2746 or 5530(2821)* 5523(1158)* ; 5532(2946)
g2747 not 2001(2825) ; 2002(2947)
g2748 or 5472(2822)* 5465(885)* ; 5474(2948)
g2749 or 4624(2829)* 4627(2827)* ; 7433(2949)
g2750 not 1751(2828) ; 1754(2950)
g2751 or 5678(2832)* 5677(2676)* ; 5679(2951)
g2752 or 5590(2833)* 5589(2677)* ; 5591(2952)
g2753 or 4989(2679)* 4988(2834)* ; 4990(2953)
g2754 or 4948(2680)* 4947(2836)* ; 4949(2954)
g2755 and 1146(2431) 1982(2816) ; 242(2955)
g2756 and 997(2432) 1790(2815) ; 266(2956)
g2757 or 3597(2841)* 3600(2838)* ; 6829(2957)
g2758 not 962(2839) ; 965(2958)
g2759 or 5108(2843)* 5107(2690)* ; 5109(2959)
g2760 or 5020(2844)* 5019(2691)* ; 5021(2960)
g2761 or 4285(2845)* 4288(2846)* ; 6337(2961)
g2762 or 1322(2847)* 1325(2848)* ; 5385(2962)
g2763 not 6362(2849) ; 6366(2963)
g2764 or 4360(2699)* 4368(2855)* ; 4381(2964)
g2765 not 6848(2851) ; 6852(2965)
g2766 and 3605(2703)* 3604(2853)* ; 3606(2966)
g2767 and 4275(2707)* 4274(2852)* ; 4276(2967)
g2768 and 4272(2710)* 4271(2857)* ; 4273(2968)
g2769 and 3602(2711)* 3601(2856)* ; 3603(2969)
g2770 and 3611(2718)* 3610(2873)* ; 3612(2970)
g2771 or 4387(2850) 4364(2720) ; 4388(2971)
g2772 and 4380(2721) 4379(2854) ; 4382(2972)
g2773 and 4638(2723)* 4637(2864)* ; 4639(2973)
g2774 or 3127(2725)* 3135(2868)* ; 3151(2974)
g2775 not 7448(2862) ; 7452(2975)
g2776 and 4635(2727)* 4634(2863)* ; 4636(2976)
g2777 and 4629(2730)* 4628(2865)* ; 4630(2977)
g2778 and 4632(2731)* 4631(2866)* ; 4633(2978)
g2779 not 6840(2867) ; 6844(2979)
g2780 or 3163(2861) 3131(2733) ; 3164(2980)
g2781 not 7458(2870) ; 7462(2981)
g2782 and 4278(2739)* 4277(2876)* ; 4279(2982)
g2783 and 4281(2740)* 4280(2872)* ; 4282(2983)
g2784 and 3608(2741)* 3607(2875)* ; 3609(2984)
g2785 not 4865(2877) ; 4871(2985)
g2786 or 6268(2808)* 6261(1944)* ; 6270(2986)
g2787 or 6179(1946)* 6176(2809)* ; 6181(2987)
g2788 or 1316(2882)* 1319(2883)* ; 5377(2988)
g2789 or 1310(2887)* 1313(2886)* ; 5369(2989)
g2790 and 3249(2223) 3035(2374) 3164(2980) ; 255(2990)
g2791 and 3249(2223) 3035(2374) 3156(2706) 4388(2971) ; 256(2991)
g2792 and 3249(2223) 3035(2374) 3164(2980) ; 261(2992)
g2793 and 3249(2223) 3035(2374) 3156(2706) 4388(2971) ; 262(2993)
g2794 not 2809(2893) ; 2812(2995)
g2795 and 4089(2553) 2854(2916) ; 1450(2996)
g2796 or 3470(2758)* 3469(2900)* ; 3471(2997)
g2797 or 3473(2759)* 3472(2901)* ; 3474(2998)
g2798 and 3466(2558) 2537(2915) ; 3274(2999)
g2799 or 3480(2765)* 3479(2902)* ; 3481(3000)
g2800 or 3477(2766)* 3476(2903)* ; 3478(3001)
g2801 or 6990(2904)* 6983(1470)* ; 6992(3002)
g2802 or 6932(2905)* 6925(1115)* ; 6934(3003)
g2803 not 3485(2909) ; 3486(3004)
g2804 not 4053(2910) ; 4056(3005)
g2805 or 7138(2913)* 7137(2780)* ; 7139(3006)
g2806 or 7050(2914)* 7049(2781)* ; 7051(3007)
g2807 and 2757(2602) 2809(2893) ; 2851(3008)
g2808 or 2542(2786)* 2541(2918)* ; 2543(3009)
g2809 or 2545(2787)* 2544(2919)* ; 2546(3010)
g2810 and 2564(2929) 2577(2920) ; 2579(3011)
g2811 or 2552(2794)* 2551(2921)* ; 2553(3012)
g2812 or 2549(2795)* 2548(2922)* ; 2550(3013)
g2813 or 6122(2923)* 6115(1494)* ; 6124(3014)
g2814 or 6064(2924)* 6057(1136)* ; 6066(3015)
g2815 and 2406(2344) 2564(2929) ; 384(3016)
g2816 not 2557(2928) ; 2558(3017)
g2817 not 2564(2929) ; 2571(3018)
g2818 not 2813(2930) ; 2816(3019)
g2819 or 4847(2932)* 4844(2345)* ; 386(3020)
g2820 or 4855(2935)* 4852(2352)* ; 389(3021)
g2821 or 4863(2938)* 4860(2358)* ; 392(3022)
g2822 or 4871(2985)* 4868(2371)* ; 395(3023)
g2823 or 7442(2814)* 7433(2949)* ; 4516(3024)
g2824 and 3035(2374) 3164(2980) ; 3239(3025)
g2825 and 3035(2374) 3156(2706) 4388(2971) ; 3240(3026)
g2826 and 997(2432) 1788(2375) 4091(2899) ; 267(3027)
g2827 and 997(2432) 1788(2375) 4089(2553) 2854(2916) ; 268(3028)
g2828 and 1788(2375) 4091(2899) ; 1436(3029)
g2829 and 1788(2375) 4089(2553) 2854(2916) ; 1440(3030)
g2830 not 1990(2943) ; 1991(3031)
g2831 and 1146(2431) 1974(2382) 3468(2898) ; 243(3032)
g2832 and 1146(2431) 1974(2382) 3466(2558) 2537(2915) ; 244(3033)
g2833 and 1974(2382) 3468(2898) ; 3265(3034)
g2834 and 1974(2382) 3466(2558) 2537(2915) ; 3267(3035)
g2835 not 1997(2944) ; 1998(3036)
g2836 or 5532(2946)* 5531(2823)* ; 5533(3037)
g2837 or 5474(2948)* 5473(2826)* ; 5475(3038)
g2838 not 7433(2949) ; 7441(3039)
g2839 or 5686(2830)* 5679(2951)* ; 5688(3040)
g2840 or 5598(2831)* 5591(2952)* ; 5600(3041)
g2841 not 5679(2951) ; 5685(3042)
g2842 not 5591(2952) ; 5597(3043)
g2843 or 6836(1833)* 6829(2957)* ; 3614(3044)
g2844 not 4990(2953) ; 4996(3045)
g2845 not 4949(2954) ; 4955(3046)
g2846 or 4997(1555)* 4990(2953)* ; 4999(3047)
g2847 or 4956(1556)* 4949(2954)* ; 4958(3048)
g2848 not 6829(2957) ; 6835(3049)
g2849 or 5116(2840)* 5109(2959)* ; 5118(3050)
g2850 or 5028(2842)* 5021(2960)* ; 5030(3051)
g2851 not 5109(2959) ; 5115(3052)
g2852 not 5021(2960) ; 5027(3053)
g2853 not 6337(2961) ; 6345(3054)
g2854 not 5385(2962) ; 5391(3055)
g2855 or 3603(2969)* 3606(2966)* ; 6837(3056)
g2856 or 4273(2968)* 4276(2967)* ; 6347(3057)
g2857 or 3609(2984)* 3612(2970)* ; 6845(3058)
g2858 and 4364(2720) 4382(2972) ; 3148(3059)
g2859 not 4382(2972) ; 4385(3060)
g2860 or 4636(2976)* 4639(2973)* ; 7443(3061)
g2861 or 4630(2977)* 4633(2978)* ; 7453(3062)
g2862 or 4279(2982)* 4282(2983)* ; 6357(3063)
g2863 or 6270(2986)* 6269(2878)* ; 6271(3064)
g2864 or 6180(2936)* 6173(1723)* ; 6182(3065)
g2865 not 5377(2988) ; 5383(3066)
g2866 or 5384(1953)* 5377(2988)* ; 1330(3067)
g2867 or 6346(2884)* 6337(2961)* ; 2860(3068)
g2868 or 5392(2885)* 5385(2962)* ; 1333(3069)
g2869 not 5369(2989) ; 5375(3070)
g2870 or 5376(1961)* 5369(2989)* ; 1327(3071)
g2871 or 3277(2891) 3274(2999) 3468(2898) ; 3279(3072)
g2872 or 1454(2894) 1450(2996) 4091(2899) ; 1766(3073)
g2873 not 3474(2998) ; 3475(3074)
g2874 not 3481(3000) ; 3482(3075)
g2875 or 6992(3002)* 6991(2907)* ; 6993(3076)
g2876 or 6934(3003)* 6933(2908)* ; 6935(3077)
g2877 or 7146(2911)* 7139(3006)* ; 7148(3078)
g2878 or 7058(2912)* 7051(3007)* ; 7060(3079)
g2879 not 7139(3006) ; 7145(3080)
g2880 not 7051(3007) ; 7057(3081)
g2881 and 2571(3018) 2495(2601) ; 2578(3082)
g2882 and 2812(2995) 2808(2917) ; 2850(3083)
g2883 not 2546(3010) ; 2547(3084)
g2884 not 2553(3012) ; 2554(3085)
g2885 and 2571(3018) 2561(2925) ; 380(3086)
g2886 or 6124(3014)* 6123(2926)* ; 6125(3087)
g2887 or 6066(3015)* 6065(2927)* ; 6067(3088)
g2888 and 2571(3018) 2400(1988) ; 383(3089)
g2889 and 2543(3009) 2564(2929) ; 375(3090)
g2890 and 2550(3013) 2564(2929) ; 378(3091)
g2891 and 2558(3017) 2564(2929) ; 381(3092)
g2892 or 6278(2940)* 6271(3064)* ; 6280(3096)
g2893 or 3241(2859) 3240(3026) 3239(3025) 3046(2813) ; 3242(3098)
g2894 or 7441(3039)* 7438(2650)* ; 4515(3099)
g2895 or 1445(2895) 1440(3030) 1436(3029) 1790(2815) ; 1447(3100)
g2896 or 3270(2892) 3267(3035) 3265(3034) 1982(2816) ; 3271(3101)
g2897 or 5540(2660)* 5533(3037)* ; 5542(3102)
g2898 or 5482(2661)* 5475(3038)* ; 5484(3103)
g2899 not 5533(3037) ; 5539(3104)
g2900 not 5475(3038) ; 5481(3105)
g2901 or 5685(3042)* 5682(2674)* ; 5687(3106)
g2902 or 5597(3043)* 5594(2675)* ; 5599(3107)
g2903 or 6835(3049)* 6832(1546)* ; 3613(3108)
g2904 or 4996(3045)* 4993(1203)* ; 4998(3111)
g2905 or 4955(3046)* 4952(1204)* ; 4957(3112)
g2906 or 5115(3052)* 5112(2687)* ; 5117(3113)
g2907 or 5027(3053)* 5024(2689)* ; 5029(3114)
g2908 or 6366(2963)* 6357(3063)* ; 2866(3115)
g2909 and 4385(3060) 4381(2964) ; 3147(3116)
g2910 or 6852(2965)* 6845(3058)* ; 3620(3117)
g2911 not 6837(3056) ; 6843(3118)
g2912 not 6347(3057) ; 6355(3119)
g2913 not 6845(3058) ; 6851(3120)
g2914 not 7443(3061) ; 7451(3123)
g2915 or 7452(2975)* 7443(3061)* ; 4519(3124)
g2916 not 7453(3062) ; 7461(3125)
g2917 or 6844(2979)* 6837(3056)* ; 3617(3126)
g2918 or 6356(2869)* 6347(3057)* ; 2863(3127)
g2919 or 7462(2981)* 7453(3062)* ; 4522(3128)
g2920 not 6357(3063) ; 6365(3129)
g2921 not 6271(3064) ; 6277(3130)
g2922 or 6182(3065)* 6181(2987)* ; 6183(3131)
g2923 or 5383(3066)* 5380(1736)* ; 1329(3132)
g2924 or 6345(3054)* 6342(2750)* ; 2859(3133)
g2925 or 5391(3055)* 5388(2751)* ; 1332(3134)
g2926 or 5375(3070)* 5372(1759)* ; 1326(3135)
g2927 and 3279(3072) ; 4713(3136)
g2928 not 1766(3073) ; 1771(3137)
g2929 or 7000(2763)* 6993(3076)* ; 7002(3138)
g2930 or 6942(2764)* 6935(3077)* ; 6944(3139)
g2931 not 6993(3076) ; 6999(3140)
g2932 not 6935(3077) ; 6941(3141)
g2933 or 7145(3080)* 7142(2778)* ; 7147(3142)
g2934 or 7057(3081)* 7054(2779)* ; 7059(3143)
g2935 or 2851(3008) 2850(3083) ; 4067(3144)
g2936 or 2579(3011) 2578(3082) ; 2580(3145)
g2937 or 6132(2792)* 6125(3087)* ; 6134(3146)
g2938 or 6074(2793)* 6067(3088)* ; 6076(3147)
g2939 not 6125(3087) ; 6131(3149)
g2940 not 6067(3088) ; 6073(3150)
g2941 and 2571(3018) 2547(3084) ; 374(3152)
g2942 and 2571(3018) 2554(3085) ; 377(3153)
g2943 or 6190(2939)* 6183(3131)* ; 6192(3154)
g2944 or 6277(3130)* 6274(2812)* ; 6279(3155)
g2945 or 4516(3024)* 4515(3099)* ; 4517(3156)
g2946 and 1447(3100) ; 975(3157)
g2947 and 3271(3101) ; 4753(3158)
g2948 or 5539(3104)* 5536(2387)* ; 5541(3159)
g2949 or 5481(3105)* 5478(2388)* ; 5483(3160)
g2950 and 3279(3072) 1950(2047) ; 2007(3161)
g2951 and 1869(1819) 1903(1826) 1885(1825) 1921(1832) 3279(3072) ; 1964(3162)
g2952 and 1903(1826) 1885(1825) 1921(1832) 3279(3072) ; 1968(3163)
g2953 or 5688(3040)* 5687(3106)* ; 5689(3164)
g2954 and 1903(1826) 1921(1832) 3279(3072) ; 1971(3165)
g2955 or 5600(3041)* 5599(3107)* ; 5601(3166)
g2956 and 1921(1832) 3279(3072) ; 1973(3167)
g2957 or 3614(3044)* 3613(3108)* ; 3615(3168)
g2958 or 4999(3047)* 4998(3111)* ; 5000(3169)
g2959 or 4958(3048)* 4957(3112)* ; 4959(3170)
g2960 or 3242(3098)* 3228(2097)* ; 3243(3171)
g2961 or 1447(3100)* 920(2100)* ; 955(3172)
g2962 and 3271(3101) 1122(2101) ; 1160(3173)
g2963 and 1038(1843) 1074(1846) 1055(1875) 1093(1853) 3271(3101) ; 1136(3174)
g2964 or 5118(3050)* 5117(3113)* ; 5119(3175)
g2965 and 1074(1846) 1055(1875) 1093(1853) 3271(3101) ; 1140(3176)
g2966 and 1074(1846) 1093(1853) 3271(3101) ; 1143(3177)
g2967 or 5030(3051)* 5029(3114)* ; 5031(3178)
g2968 and 1093(1853) 3271(3101) ; 1145(3179)
g2969 or 6365(3129)* 6362(2849)* ; 2865(3180)
g2970 or 6851(3120)* 6848(2851)* ; 3619(3181)
g2971 or 3148(3059) 3147(3116) ; 3149(3182)
g2972 or 7451(3123)* 7448(2862)* ; 4518(3183)
g2973 or 6843(3118)* 6840(2867)* ; 3616(3184)
g2974 or 6355(3119)* 6352(2734)* ; 2862(3185)
g2975 or 7461(3125)* 7458(2870)* ; 4521(3186)
g2976 not 6183(3131) ; 6189(3187)
g2977 or 1330(3067)* 1329(3132)* ; 1331(3188)
g2978 or 2860(3068)* 2859(3133)* ; 2861(3189)
g2979 or 1333(3069)* 1332(3134)* ; 1334(3190)
g2980 or 1327(3071)* 1326(3135)* ; 1328(3191)
g2981 not 4713(3136) ; 4719(3192)
g2982 or 6999(3140)* 6996(2561)* ; 7001(3193)
g2983 or 6941(3141)* 6938(2562)* ; 6943(3194)
g2984 and 2580(3145) 3446(2265) ; 3490(3195)
g2985 and 3365(1973) 3399(1978) 3381(1976) 3417(1979) 2580(3145) ; 3459(3196)
g2986 and 3399(1978) 3381(1976) 3417(1979) 2580(3145) ; 3462(3197)
g2987 or 7148(3078)* 7147(3142)* ; 7149(3198)
g2988 or 7060(3079)* 7059(3143)* ; 7061(3199)
g2989 and 3399(1978) 3417(1979) 2580(3145) ; 3464(3200)
g2990 and 3417(1979) 2580(3145) ; 3465(3201)
g2991 not 4067(3144) ; 4072(3202)
g2992 and 2580(3145) ; 4793(3203)
g2993 or 6131(3149)* 6128(2611)* ; 6133(3204)
g2994 or 6073(3150)* 6070(2612)* ; 6075(3205)
g2995 or 6189(3187)* 6186(2811)* ; 6191(3208)
g2996 or 6280(3096)* 6279(3155)* ; 6281(3209)
g2997 not 975(3157) ; 980(3210)
g2998 not 4753(3158) ; 4759(3211)
g2999 or 5542(3102)* 5541(3159)* ; 5543(3212)
g3000 or 5484(3103)* 5483(3160)* ; 5485(3213)
g3001 or 2007(3161) 1957(2411) ; 2008(3214)
g3002 or 5696(2669)* 5689(3164)* ; 5698(3215)
g3003 or 5608(2670)* 5601(3166)* ; 5610(3216)
g3004 or 1964(3162) 1962(2086) 1961(2072) 1960(2059) 1880(895) ; 4721(3217)
g3005 or 1968(3163) 1966(2089) 1965(2074) 1897(900) ; 4729(3218)
g3006 not 5689(3164) ; 5695(3219)
g3007 or 1971(3165) 1969(2088) 1914(905) ; 4737(3220)
g3008 not 5601(3166) ; 5607(3221)
g3009 or 1973(3167) 1929(910) ; 4745(3222)
g3010 or 4720(2430)* 4713(3136)* ; 294(3223)
g3011 or 4966(1198)* 4959(3170)* ; 4968(3224)
g3012 or 5007(1201)* 5000(3169)* ; 5009(3225)
g3013 not 5000(3169) ; 5006(3226)
g3014 not 4959(3170) ; 4965(3227)
g3015 and 955(3172) 933(2683) ; 958(3228)
g3016 or 1160(3173) 1129(2434) ; 1161(3229)
g3017 and 3243(3171) 3238(2684) ; 3245(3230)
g3018 or 5126(2685)* 5119(3175)* ; 5128(3231)
g3019 or 5038(2686)* 5031(3178)* ; 5040(3232)
g3020 or 1136(3174) 1134(2131) 1133(2115) 1132(2164) 1050(930) ; 4761(3233)
g3021 not 5119(3175) ; 5125(3234)
g3022 or 1143(3177) 1141(2133) 1086(935) ; 4777(3235)
g3023 not 5031(3178) ; 5037(3236)
g3024 or 1145(3179) 1102(940) ; 4785(3237)
g3025 or 4760(2455)* 4753(3158)* ; 323(3238)
g3026 or 2866(3115)* 2865(3180)* ; 2867(3239)
g3027 or 3620(3117)* 3619(3181)* ; 3621(3240)
g3028 or 3149(3182)* 3136(2475)* ; 3150(3241)
g3029 or 1140(3176) 1138(2134) 1137(2117) 1068(981) ; 4769(3242)
g3030 or 4519(3124)* 4518(3183)* ; 4520(3243)
g3031 or 3617(3126)* 3616(3184)* ; 3618(3244)
g3032 or 2863(3127)* 2862(3185)* ; 2864(3245)
g3033 or 4522(3128)* 4521(3186)* ; 4523(3246)
g3034 or 7002(3138)* 7001(3193)* ; 7003(3247)
g3035 or 6944(3139)* 6943(3194)* ; 6945(3248)
g3036 or 3490(3195) 3453(2578) ; 3491(3249)
g3037 or 3459(3196) 3458(2294) 3457(2282) 3456(2273) 3376(1119) ; 4801(3250)
g3038 or 7156(2774)* 7149(3198)* ; 7158(3251)
g3039 or 7068(2775)* 7061(3199)* ; 7070(3252)
g3040 or 3462(3197) 3461(2297) 3460(2284) 3393(1121) ; 4809(3253)
g3041 or 3464(3200) 3463(2296) 3410(1123) ; 4817(3254)
g3042 not 7149(3198) ; 7155(3255)
g3043 not 7061(3199) ; 7067(3256)
g3044 or 3465(3201) 3425(1125) ; 4825(3257)
g3045 or 4800(2598)* 4793(3203)* ; 343(3258)
g3046 not 4793(3203) ; 4799(3259)
g3047 or 6134(3146)* 6133(3204)* ; 6135(3260)
g3048 or 6076(3147)* 6075(3205)* ; 6077(3261)
g3049 or 6288(2805)* 6281(3209)* ; 6290(3262)
g3050 or 6192(3154)* 6191(3208)* ; 6193(3263)
g3051 not 6281(3209) ; 6287(3264)
g3052 and 4523(3246) 4520(3243) 4517(3156) 3615(3168) ; 4524(3265)
g3053 and 1987(2942) 2008(3214) ; 297(3266)
g3054 and 1994(2945) 2008(3214) ; 300(3267)
g3055 not 5543(3212) ; 5549(3268)
g3056 not 5485(3213) ; 5491(3269)
g3057 and 1856(2037) 2008(3214) ; 306(3270)
g3058 and 2002(2947) 2008(3214) ; 303(3271)
g3059 or 5550(2401)* 5543(3212)* ; 5552(3272)
g3060 or 5492(2402)* 5485(3213)* ; 5494(3273)
g3061 not 2008(3214) ; 2014(3274)
g3062 or 4728(2412)* 4721(3217)* ; 309(3275)
g3063 or 5695(3219)* 5692(2413)* ; 5697(3276)
g3064 or 5607(3221)* 5604(2414)* ; 5609(3277)
g3065 not 4721(3217) ; 4727(3278)
g3066 or 4736(2415)* 4729(3218)* ; 312(3279)
g3067 not 4729(3218) ; 4735(3280)
g3068 or 4744(2423)* 4737(3220)* ; 315(3281)
g3069 not 4737(3220) ; 4743(3282)
g3070 or 4752(2425)* 4745(3222)* ; 318(3283)
g3071 not 4745(3222) ; 4751(3284)
g3072 or 4719(3192)* 4716(2094)* ; 293(3285)
g3073 and 908(1192) 958(3228) ; 275(3286)
g3074 and 1161(3229) 1176(1838) ; 272(3287)
g3075 or 4965(3227)* 4962(919)* ; 4967(3288)
g3076 or 5006(3226)* 5003(920)* ; 5008(3289)
g3077 and 1023(1205) 1161(3229) ; 1174(3290)
g3078 not 958(3228) ; 961(3291)
g3079 not 1161(3229) ; 1166(3292)
g3080 not 3245(3230) ; 3248(3293)
g3081 or 4768(2442)* 4761(3233)* ; 326(3294)
g3082 or 5125(3234)* 5122(2443)* ; 5127(3295)
g3083 or 5037(3236)* 5034(2444)* ; 5039(3296)
g3084 not 4761(3233) ; 4767(3297)
g3085 or 4776(2445)* 4769(3242)* ; 329(3298)
g3086 not 4777(3235) ; 4783(3299)
g3087 or 4792(2449)* 4785(3237)* ; 335(3300)
g3088 not 4785(3237) ; 4791(3301)
g3089 or 4759(3211)* 4756(2139)* ; 322(3302)
g3090 not 4769(3242) ; 4775(3303)
g3091 or 4784(2485)* 4777(3235)* ; 332(3304)
g3092 and 3150(3241) 3146(2871) ; 3152(3305)
g3093 and 3223(1698) 3245(3230) ; 248(3306)
g3094 and 1155(2201) 1161(3229) ; 1171(3307)
g3095 and 2867(3239) 2864(3245) 2861(3189) 1331(3188) ; 2868(3308)
g3096 and 3621(3240) 3618(3244) 1334(3190) 1328(3191) ; 4443(3309)
g3097 and 3248(3293) 3244(1962) ; 247(3310)
g3098 and 3471(2997) 3491(3249) ; 346(3311)
g3099 not 7003(3247) ; 7009(3312)
g3100 not 6945(3248) ; 6951(3313)
g3101 and 3478(3001) 3491(3249) ; 349(3314)
g3102 or 7010(2575)* 7003(3247)* ; 7012(3315)
g3103 or 6952(2576)* 6945(3248)* ; 6954(3316)
g3104 and 3350(2261) 3491(3249) ; 355(3317)
g3105 and 3486(3004) 3491(3249) ; 352(3318)
g3106 not 3491(3249) ; 3497(3319)
g3107 or 4808(2583)* 4801(3250)* ; 358(3320)
g3108 not 4801(3250) ; 4807(3321)
g3109 or 7155(3255)* 7152(2584)* ; 7157(3322)
g3110 or 7067(3256)* 7064(2585)* ; 7069(3323)
g3111 or 4816(2586)* 4809(3253)* ; 361(3324)
g3112 not 4809(3253) ; 4815(3325)
g3113 or 4824(2593)* 4817(3254)* ; 364(3326)
g3114 not 4817(3254) ; 4823(3327)
g3115 or 4832(2597)* 4825(3257)* ; 367(3328)
g3116 not 4825(3257) ; 4831(3329)
g3117 or 4799(3259)* 4796(2304)* ; 342(3330)
g3118 not 6135(3260) ; 6141(3331)
g3119 not 6077(3261) ; 6083(3332)
g3120 or 6142(2625)* 6135(3260)* ; 6144(3333)
g3121 or 6084(2626)* 6077(3261)* ; 6086(3334)
g3122 or 6287(3264)* 6284(2635)* ; 6289(3335)
g3123 or 6200(2933)* 6193(3263)* ; 6202(3336)
g3124 not 6193(3263) ; 6199(3337)
g3125 and 2868(3308) 4524(3265) 4443(3309) ; 2881(3339)
g3126 and 2014(3274) 1991(3031) ; 296(3340)
g3127 and 2014(3274) 1998(3036) ; 299(3341)
g3128 and 2014(3274) 2005(2824) ; 302(3342)
g3129 and 2014(3274) 1850(1812) ; 305(3343)
g3130 or 5549(3268)* 5546(2038)* ; 5551(3344)
g3131 or 5491(3269)* 5488(2039)* ; 5493(3345)
g3132 or 4727(3278)* 4724(2048)* ; 308(3346)
g3133 or 5698(3215)* 5697(3276)* ; 5699(3347)
g3134 or 5610(3216)* 5609(3277)* ; 5611(3348)
g3135 or 4735(3280)* 4732(2051)* ; 311(3349)
g3136 or 4743(3282)* 4740(2066)* ; 314(3350)
g3137 or 4751(3284)* 4748(2075)* ; 317(3351)
g3138 and 961(3291) 957(1836) ; 274(3353)
g3139 and 1166(3292) 1117(1193) ; 271(3354)
g3140 or 4968(3224)* 4967(3288)* ; 967(3355)
g3141 or 5009(3225)* 5008(3289)* ; 971(3356)
g3142 and 1166(3292) 1019(923) ; 1173(3357)
g3143 or 4767(3297)* 4764(2102)* ; 325(3358)
g3144 or 5128(3231)* 5127(3295)* ; 5129(3359)
g3145 or 5040(3232)* 5039(3296)* ; 5041(3360)
g3146 or 4775(3303)* 4772(2105)* ; 328(3361)
g3147 or 4791(3301)* 4788(2118)* ; 334(3362)
g3148 or 4783(3299)* 4780(2168)* ; 331(3364)
g3149 and 3131(2733) 3152(3305) ; 251(3365)
g3150 not 3152(3305) ; 3155(3366)
g3151 and 1166(3292) 1158(1927) ; 1170(3367)
g3152 and 3497(3319) 3475(3074) ; 345(3370)
g3153 and 3497(3319) 3482(3075) ; 348(3371)
g3154 and 3497(3319) 3489(2906) ; 351(3372)
g3155 or 7009(3312)* 7006(2259)* ; 7011(3373)
g3156 or 6951(3313)* 6948(2260)* ; 6953(3374)
g3157 and 3497(3319) 3344(1970) ; 354(3375)
g3158 or 4807(3321)* 4804(2266)* ; 357(3376)
g3159 or 7158(3251)* 7157(3322)* ; 7159(3377)
g3160 or 7070(3252)* 7069(3323)* ; 7071(3378)
g3161 or 4815(3325)* 4812(2269)* ; 360(3379)
g3162 or 4823(3327)* 4820(2281)* ; 363(3380)
g3163 or 4831(3329)* 4828(2293)* ; 366(3381)
g3164 or 6141(3331)* 6138(2342)* ; 6143(3383)
g3165 or 6083(3332)* 6080(2343)* ; 6085(3384)
g3166 or 6290(3262)* 6289(3335)* ; 6291(3385)
g3167 or 6199(3337)* 6196(2806)* ; 6201(3386)
g3168 or 5552(3272)* 5551(3344)* ; 5553(3391)
g3169 or 5494(3273)* 5493(3345)* ; 5495(3392)
g3170 not 5699(3347) ; 5705(3394)
g3171 not 5611(3348) ; 5617(3395)
g3172 or 5706(2428)* 5699(3347)* ; 5708(3399)
g3173 or 5618(2429)* 5611(3348)* ; 5620(3400)
g3174 or 1174(3290) 1173(3357) ; 1175(3403)
g3175 and 980(3210) 929(2433) 967(3355) ; 992(3404)
g3176 and 980(3210) 933(2683) 971(3356) ; 991(3405)
g3177 and 975(3157) 962(2839) 971(3356) ; 993(3406)
g3178 and 975(3157) 965(2958) 967(3355) ; 994(3407)
g3179 not 5129(3359) ; 5135(3409)
g3180 not 5041(3360) ; 5047(3410)
g3181 or 5136(2453)* 5129(3359)* ; 5138(3413)
g3182 or 5048(2454)* 5041(3360)* ; 5050(3414)
g3183 and 2881(3339) 2878(386) 2876(389) ; 417(3415)
g3184 and 3155(3366) 3151(2974) ; 250(3417)
g3185 or 1171(3307) 1170(3367) ; 1172(3419)
g3186 or 7012(3315)* 7011(3373)* ; 7013(3422)
g3187 or 6954(3316)* 6953(3374)* ; 6955(3423)
g3188 not 7159(3377) ; 7165(3427)
g3189 not 7071(3378) ; 7077(3428)
g3190 or 7166(2599)* 7159(3377)* ; 7168(3432)
g3191 or 7078(2600)* 7071(3378)* ; 7080(3433)
g3192 or 6144(3333)* 6143(3383)* ; 6145(3434)
g3193 or 6086(3334)* 6085(3384)* ; 6087(3435)
g3194 not 6291(3385) ; 6297(3436)
g3195 or 6202(3336)* 6201(3386)* ; 6203(3437)
g3196 or 5502(2395)* 5495(3392)* ; 5504(3438)
g3197 or 5560(2396)* 5553(3391)* ; 5562(3439)
g3198 not 5553(3391) ; 5559(3440)
g3199 not 5495(3392) ; 5501(3441)
g3200 or 5705(3394)* 5702(2090)* ; 5707(3442)
g3201 or 5617(3395)* 5614(2091)* ; 5619(3443)
g3202 or 994(3407) 993(3406) 992(3404) 991(3405) ; 5167(3446)
g3203 or 5135(3409)* 5132(2135)* ; 5137(3447)
g3204 or 5047(3410)* 5044(2136)* ; 5049(3448)
g3205 or 6298(2880)* 6291(3385)* ; 6300(3453)
g3206 or 6962(2572)* 6955(3423)* ; 6964(3454)
g3207 or 7020(2573)* 7013(3422)* ; 7022(3455)
g3208 not 7013(3422) ; 7019(3456)
g3209 not 6955(3423) ; 6961(3457)
g3210 or 7165(3427)* 7162(2305)* ; 7167(3458)
g3211 or 7077(3428)* 7074(2306)* ; 7079(3459)
g3212 or 6094(2620)* 6087(3435)* ; 6096(3460)
g3213 or 6152(2621)* 6145(3434)* ; 6154(3461)
g3214 not 6145(3434) ; 6151(3462)
g3215 not 6087(3435) ; 6093(3463)
g3216 not 6203(3437) ; 6209(3464)
g3217 or 5501(3441)* 5498(2023)* ; 5503(3465)
g3218 or 5559(3440)* 5556(2024)* ; 5561(3466)
g3219 or 5708(3399)* 5707(3442)* ; 5709(3467)
g3220 or 5620(3400)* 5619(3443)* ; 5621(3468)
g3221 not 5167(3446) ; 5173(3469)
g3222 or 5138(3413)* 5137(3447)* ; 5139(3470)
g3223 or 5050(3414)* 5049(3448)* ; 5051(3471)
g3224 or 6297(3436)* 6294(2746)* ; 6299(3472)
g3225 or 6210(2881)* 6203(3437)* ; 6212(3473)
g3226 or 6961(3457)* 6958(2248)* ; 6963(3474)
g3227 or 7019(3456)* 7016(2249)* ; 7021(3475)
g3228 or 7168(3432)* 7167(3458)* ; 7169(3476)
g3229 or 7080(3433)* 7079(3459)* ; 7081(3477)
g3230 or 6093(3463)* 6090(2328)* ; 6095(3478)
g3231 or 6151(3462)* 6148(2329)* ; 6153(3479)
g3232 or 5504(3438)* 5503(3465)* ; 5505(3480)
g3233 or 5562(3439)* 5561(3466)* ; 5563(3481)
g3234 or 5628(2426)* 5621(3468)* ; 5630(3482)
g3235 or 5716(2427)* 5709(3467)* ; 5718(3483)
g3236 not 5709(3467) ; 5715(3484)
g3237 not 5621(3468) ; 5627(3485)
g3238 or 5058(2451)* 5051(3471)* ; 5060(3486)
g3239 or 5146(2452)* 5139(3470)* ; 5148(3487)
g3240 not 5139(3470) ; 5145(3488)
g3241 not 5051(3471) ; 5057(3489)
g3242 or 6300(3453)* 6299(3472)* ; 6301(3490)
g3243 or 6209(3464)* 6206(2747)* ; 6211(3491)
g3244 or 6964(3454)* 6963(3474)* ; 6965(3492)
g3245 or 7022(3455)* 7021(3475)* ; 7023(3493)
g3246 or 7088(2595)* 7081(3477)* ; 7090(3494)
g3247 or 7176(2596)* 7169(3476)* ; 7178(3495)
g3248 not 7169(3476) ; 7175(3496)
g3249 not 7081(3477) ; 7087(3497)
g3250 or 6096(3460)* 6095(3478)* ; 6097(3498)
g3251 or 6154(3461)* 6153(3479)* ; 6155(3499)
g3252 or 6308(2647)* 6301(3490)* ; 6310(3500)
g3253 or 5570(2376)* 5563(3481)* ; 5572(3501)
g3254 or 5512(2377)* 5505(3480)* ; 5514(3502)
g3255 not 5505(3480) ; 5511(3503)
g3256 not 5563(3481) ; 5569(3504)
g3257 or 5627(3485)* 5624(2076)* ; 5629(3505)
g3258 or 5715(3484)* 5712(2077)* ; 5717(3506)
g3259 or 5057(3489)* 5054(2121)* ; 5059(3507)
g3260 or 5145(3488)* 5142(2123)* ; 5147(3508)
g3261 not 6301(3490) ; 6307(3509)
g3262 or 6212(3473)* 6211(3491)* ; 6213(3510)
g3263 or 7030(2554)* 7023(3493)* ; 7032(3511)
g3264 or 6972(2555)* 6965(3492)* ; 6974(3512)
g3265 not 6965(3492) ; 6971(3513)
g3266 not 7023(3493) ; 7029(3514)
g3267 or 7087(3497)* 7084(2290)* ; 7089(3515)
g3268 or 7175(3496)* 7172(2291)* ; 7177(3516)
g3269 or 6162(2604)* 6155(3499)* ; 6164(3517)
g3270 or 6104(2605)* 6097(3498)* ; 6106(3518)
g3271 not 6097(3498) ; 6103(3519)
g3272 not 6155(3499) ; 6161(3520)
g3273 or 6220(2646)* 6213(3510)* ; 6222(3521)
g3274 or 6307(3509)* 6304(2370)* ; 6309(3522)
g3275 or 5569(3504)* 5566(2000)* ; 5571(3523)
g3276 or 5511(3503)* 5508(2001)* ; 5513(3524)
g3277 or 5630(3482)* 5629(3505)* ; 5631(3525)
g3278 or 5718(3483)* 5717(3506)* ; 5719(3526)
g3279 or 5060(3486)* 5059(3507)* ; 5061(3527)
g3280 or 5148(3487)* 5147(3508)* ; 5149(3528)
g3281 not 6213(3510) ; 6219(3529)
g3282 or 7029(3514)* 7026(2225)* ; 7031(3530)
g3283 or 6971(3513)* 6968(2226)* ; 6973(3531)
g3284 or 7090(3494)* 7089(3515)* ; 7091(3532)
g3285 or 7178(3495)* 7177(3516)* ; 7179(3533)
g3286 or 6161(3520)* 6158(2308)* ; 6163(3534)
g3287 or 6103(3519)* 6100(2309)* ; 6105(3535)
g3288 or 6219(3529)* 6216(2369)* ; 6221(3536)
g3289 or 6310(3500)* 6309(3522)* ; 6311(3537)
g3290 or 5572(3501)* 5571(3523)* ; 5573(3538)
g3291 or 5514(3502)* 5513(3524)* ; 5515(3539)
g3292 or 5726(2408)* 5719(3526)* ; 5728(3540)
g3293 or 5638(2409)* 5631(3525)* ; 5640(3541)
g3294 not 5631(3525) ; 5637(3542)
g3295 not 5719(3526) ; 5725(3543)
g3296 or 5156(2439)* 5149(3528)* ; 5158(3544)
g3297 or 5068(2440)* 5061(3527)* ; 5070(3545)
g3298 not 5061(3527) ; 5067(3546)
g3299 not 5149(3528) ; 5155(3547)
g3300 or 7032(3511)* 7031(3530)* ; 7033(3548)
g3301 or 6974(3512)* 6973(3531)* ; 6975(3549)
g3302 or 7186(2580)* 7179(3533)* ; 7188(3550)
g3303 or 7098(2581)* 7091(3532)* ; 7100(3551)
g3304 not 7091(3532) ; 7097(3552)
g3305 not 7179(3533) ; 7185(3553)
g3306 or 6164(3517)* 6163(3534)* ; 6165(3554)
g3307 or 6106(3518)* 6105(3535)* ; 6107(3555)
g3308 or 6318(2632)* 6311(3537)* ; 6320(3556)
g3309 or 6222(3521)* 6221(3536)* ; 6223(3557)
g3310 not 6311(3537) ; 6317(3558)
g3311 not 5573(3538) ; 5579(3559)
g3312 not 5515(3539) ; 5521(3560)
g3313 or 5522(2389)* 5515(3539)* ; 1756(3561)
g3314 or 5580(2390)* 5573(3538)* ; 1761(3562)
g3315 or 5725(3543)* 5722(2044)* ; 5727(3563)
g3316 or 5637(3542)* 5634(2045)* ; 5639(3564)
g3317 or 5155(3547)* 5152(2098)* ; 5157(3565)
g3318 or 5067(3546)* 5064(2099)* ; 5069(3566)
g3319 not 7033(3548) ; 7039(3567)
g3320 not 6975(3549) ; 6981(3568)
g3321 or 6982(2565)* 6975(3549)* ; 4058(3569)
g3322 or 7040(2566)* 7033(3548)* ; 4063(3570)
g3323 or 7185(3553)* 7182(2262)* ; 7187(3571)
g3324 or 7097(3552)* 7094(2263)* ; 7099(3572)
g3325 not 6165(3554) ; 6171(3573)
g3326 not 6107(3555) ; 6113(3574)
g3327 or 6114(2615)* 6107(3555)* ; 2818(3575)
g3328 or 6172(2616)* 6165(3554)* ; 2823(3576)
g3329 or 6317(3558)* 6314(2346)* ; 6319(3577)
g3330 or 6230(2633)* 6223(3557)* ; 6232(3578)
g3331 not 6223(3557) ; 6229(3579)
g3332 or 5521(3560)* 5518(2011)* ; 1755(3580)
g3333 or 5579(3559)* 5576(2013)* ; 1760(3581)
g3334 or 5728(3540)* 5727(3563)* ; 5729(3582)
g3335 or 5640(3541)* 5639(3564)* ; 5641(3583)
g3336 or 5158(3544)* 5157(3565)* ; 5159(3584)
g3337 or 5070(3545)* 5069(3566)* ; 5071(3585)
g3338 or 6981(3568)* 6978(2235)* ; 4057(3586)
g3339 or 7039(3567)* 7036(2237)* ; 4062(3587)
g3340 or 7188(3550)* 7187(3571)* ; 7189(3588)
g3341 or 7100(3551)* 7099(3572)* ; 7101(3589)
g3342 or 6113(3574)* 6110(2318)* ; 2817(3590)
g3343 or 6171(3573)* 6168(2320)* ; 2822(3591)
g3344 or 6320(3556)* 6319(3577)* ; 6321(3592)
g3345 or 6229(3579)* 6226(2347)* ; 6231(3593)
g3346 or 1756(3561)* 1755(3580)* ; 1757(3594)
g3347 or 1761(3562)* 1760(3581)* ; 1762(3595)
g3348 not 5729(3582) ; 5735(3596)
g3349 not 5641(3583) ; 5647(3597)
g3350 or 5736(2421)* 5729(3582)* ; 5660(3598)
g3351 or 5648(2422)* 5641(3583)* ; 5650(3599)
g3352 not 5159(3584) ; 5165(3600)
g3353 not 5071(3585) ; 5077(3601)
g3354 or 5166(2483)* 5159(3584)* ; 5090(3602)
g3355 or 5078(2484)* 5071(3585)* ; 5080(3603)
g3356 or 4058(3569)* 4057(3586)* ; 4059(3604)
g3357 or 4063(3570)* 4062(3587)* ; 4064(3605)
g3358 not 7189(3588) ; 7195(3606)
g3359 not 7101(3589) ; 7107(3607)
g3360 or 7196(2591)* 7189(3588)* ; 7120(3608)
g3361 or 7108(2592)* 7101(3589)* ; 7110(3609)
g3362 or 2818(3575)* 2817(3590)* ; 2819(3610)
g3363 or 2823(3576)* 2822(3591)* ; 2824(3611)
g3364 not 6321(3592) ; 6327(3612)
g3365 or 6232(3578)* 6231(3593)* ; 6233(3613)
g3366 or 6328(2642)* 6321(3592)* ; 6252(3614)
g3367 and 1771(3137) 1726(2407) 1757(3594) ; 1783(3615)
g3368 and 1771(3137) 1730(2668) 1762(3595) ; 1782(3616)
g3369 and 1766(3073) 1751(2828) 1762(3595) ; 1784(3617)
g3370 and 1766(3073) 1754(2950) 1757(3594) ; 1785(3618)
g3371 or 5735(3596)* 5732(2063)* ; 5659(3619)
g3372 or 5647(3597)* 5644(2064)* ; 5649(3620)
g3373 or 5165(3600)* 5162(2166)* ; 5089(3621)
g3374 or 5077(3601)* 5074(2167)* ; 5079(3622)
g3375 and 2828(208) 2813(2930) 2824(3611) ; 2846(3623)
g3376 and 2828(208) 2816(3019) 2819(3610) ; 2847(3624)
g3377 and 2833(317) 2784(2802) 2824(3611) ; 2844(3625)
g3378 and 2833(317) 2780(2629) 2819(3610) ; 2845(3626)
g3379 and 4072(3202) 4028(2579) 4059(3604) ; 4084(3627)
g3380 and 4072(3202) 4032(2773) 4064(3605) ; 4083(3628)
g3381 and 4067(3144) 4053(2910) 4064(3605) ; 4085(3629)
g3382 and 4067(3144) 4056(3005) 4059(3604) ; 4086(3630)
g3383 or 7195(3606)* 7192(2278)* ; 7119(3631)
g3384 or 7107(3607)* 7104(2279)* ; 7109(3632)
g3385 not 6233(3613) ; 6239(3633)
g3386 or 6327(3612)* 6324(2359)* ; 6251(3634)
g3387 or 6240(2643)* 6233(3613)* ; 6242(3635)
g3388 or 1785(3618) 1784(3617) 1783(3615) 1782(3616) ; 5737(3636)
g3389 or 5660(3598)* 5659(3619)* ; 5661(3637)
g3390 or 5650(3599)* 5649(3620)* ; 5651(3638)
g3391 or 5090(3602)* 5089(3621)* ; 5091(3639)
g3392 or 5080(3603)* 5079(3622)* ; 5081(3640)
g3393 or 2847(3624) 2846(3623) 2845(3626) 2844(3625) ; 6329(3641)
g3394 or 4086(3630) 4085(3629) 4084(3627) 4083(3628) ; 7197(3642)
g3395 or 7120(3608)* 7119(3631)* ; 7121(3643)
g3396 or 7110(3609)* 7109(3632)* ; 7111(3644)
g3397 or 6252(3614)* 6251(3634)* ; 6253(3645)
g3398 or 6239(3633)* 6236(2360)* ; 6241(3646)
g3399 not 5737(3636) ; 5743(3647)
g3400 or 5668(2416)* 5661(3637)* ; 1779(3648)
g3401 or 5658(2417)* 5651(3638)* ; 1776(3649)
g3402 not 5661(3637) ; 5667(3650)
g3403 not 5651(3638) ; 5657(3651)
g3404 or 5098(2446)* 5091(3639)* ; 988(3652)
g3405 or 5088(2447)* 5081(3640)* ; 985(3653)
g3406 not 5091(3639) ; 5097(3654)
g3407 not 5081(3640) ; 5087(3655)
g3408 not 6329(3641) ; 6335(3656)
g3409 not 7197(3642) ; 7203(3657)
g3410 or 7128(2587)* 7121(3643)* ; 4080(3658)
g3411 or 7118(2588)* 7111(3644)* ; 4077(3659)
g3412 not 7121(3643) ; 7127(3660)
g3413 not 7111(3644) ; 7117(3661)
g3414 or 6260(2636)* 6253(3645)* ; 2841(3662)
g3415 not 6253(3645) ; 6259(3663)
g3416 or 6242(3635)* 6241(3646)* ; 6243(3664)
g3417 or 5667(3650)* 5664(2052)* ; 1778(3665)
g3418 or 5657(3651)* 5654(2054)* ; 1775(3666)
g3419 or 5097(3654)* 5094(2106)* ; 987(3667)
g3420 or 5087(3655)* 5084(2108)* ; 984(3668)
g3421 or 7127(3660)* 7124(2270)* ; 4079(3669)
g3422 or 7117(3661)* 7114(2272)* ; 4076(3670)
g3423 or 6259(3663)* 6256(2350)* ; 2840(3671)
g3424 or 6250(2638)* 6243(3664)* ; 2838(3672)
g3425 not 6243(3664) ; 6249(3673)
g3426 or 1779(3648)* 1778(3665)* ; 1780(3674)
g3427 or 1776(3649)* 1775(3666)* ; 1777(3675)
g3428 or 988(3652)* 987(3667)* ; 989(3676)
g3429 or 985(3653)* 984(3668)* ; 986(3677)
g3430 and 1777(3675) 1766(3073) ; 1787(3678)
g3431 or 4080(3658)* 4079(3669)* ; 4081(3679)
g3432 or 4077(3659)* 4076(3670)* ; 4078(3680)
g3433 or 2841(3662)* 2840(3671)* ; 2842(3681)
g3434 or 6249(3673)* 6246(2351)* ; 2837(3682)
g3435 and 986(3677) 975(3157) ; 996(3683)
g3436 not 1780(3674) ; 1781(3684)
g3437 not 989(3676) ; 990(3685)
g3438 and 1771(3137) 1781(3684) ; 1786(3686)
g3439 not 4081(3679) ; 4082(3687)
g3440 and 4078(3680) 4067(3144) ; 4088(3688)
g3441 not 2842(3681) ; 2843(3689)
g3442 or 2838(3672)* 2837(3682)* ; 2839(3690)
g3443 and 980(3210) 990(3685) ; 995(3691)
g3444 and 2839(3690) 2828(208) ; 2849(3692)
g3445 and 2833(317) 2843(3689) ; 2848(3693)
g3446 or 1787(3678) 1786(3686) ; 5740(3694)
g3447 and 4072(3202) 4082(3687) ; 4087(3695)
g3448 or 996(3683) 995(3691) ; 5170(3696)
g3449 or 2849(3692) 2848(3693) ; 6332(3697)
g3450 not 5740(3694) ; 5744(3698)
g3451 or 4088(3688) 4087(3695) ; 7200(3699)
g3452 not 5170(3696) ; 5174(3700)
g3453 or 5743(3647)* 5740(3694)* ; 1791(3701)
g3454 or 5173(3469)* 5170(3696)* ; 1003(3702)
g3455 or 6335(3656)* 6332(3697)* ; 2855(3703)
g3456 not 6332(3697) ; 6336(3704)
g3457 or 7203(3657)* 7200(3699)* ; 4092(3705)
g3458 not 7200(3699) ; 7204(3706)
g3459 or 5744(3698)* 5737(3636)* ; 1792(3707)
g3460 or 5174(3700)* 5167(3446)* ; 1004(3708)
g3461 or 6336(3704)* 6329(3641)* ; 2856(3709)
g3462 or 7204(3706)* 7197(3642)* ; 4093(3710)
g3463 or 1792(3707)* 1791(3701)* ; 320(3711)
g3464 or 1004(3708)* 1003(3702)* ; 337(3712)
g3465 or 2856(3709)* 2855(3703)* ; 398(3713)
g3466 or 4093(3710)* 4092(3705)* ; 369(3714)
g3467 and IN-339(164) ; 339(164)
g3468 and 1(0) ; 2(313)
g3469 and 1(0) ; 3(312)
g3470 and 1459(167) ; 450(288)
g3471 and 1469(169) ; 448(284)
g3472 and 1480(170) ; 444(282)
g3473 and 1486(171) ; 442(280)
g3474 and 1492(172) ; 440(277)
g3475 and 1496(173) ; 438(274)
g3476 and 2208(175) ; 496(271)
g3477 and 2218(177) ; 494(267)
g3478 and 2224(178) ; 492(265)
g3479 and 2230(179) ; 490(263)
g3480 and 2236(180) ; 488(260)
g3481 and 2239(181) ; 486(258)
g3482 and 2247(182) ; 484(256)
g3483 and 2253(183) ; 482(253)
g3484 and 2256(184) ; 480(250)
g3485 and 3698(185) ; 560(248)
g3486 and 3701(186) ; 542(246)
g3487 and 3705(187) ; 558(244)
g3488 and 3711(188) ; 556(242)
g3489 and 3717(189) ; 554(240)
g3490 and 3723(190) ; 552(238)
g3491 and 3729(191) ; 550(236)
g3492 and 3737(192) ; 548(234)
g3493 and 3743(193) ; 546(232)
g3494 and 3749(194) ; 544(230)
g3495 and 4393(195) ; 540(227)
g3496 and 4400(197) ; 538(224)
g3497 and 4405(198) ; 536(222)
g3498 and 4410(199) ; 534(220)
g3499 and 4415(200) ; 532(218)
g3500 and 4420(201) ; 530(216)
g3501 and 4427(202) ; 528(214)
g3502 and 4432(203) ; 526(212)
g3503 and 4437(204) ; 524(210)
g3504 and 1462(168) ; 436(286)
g3505 and 2211(176) ; 478(269)
g3506 and 4394(196) ; 522(226)
g3507 and 1172(3419) ; 422(3451)
g3508 and 1172(3419) ; 469(3452)
g3509 and 1175(3403) ; 419(3444)
g3510 and 1175(3403) ; 471(3445)
g3511 not 400(297) ; 400(297)*
g3512 not 401(310) ; 401(310)*
g3513 not 1197(165) ; 1197(165)*
g3514 not 574(308) ; 574(308)*
g3515 not 1184(294) ; 1184(294)*
g3516 not 575(309) ; 575(309)*
g3517 not 371(2754) ; 371(2754)*
g3518 not 372(2890) ; 372(2890)*
g3519 not 386(3020) ; 386(3020)*
g3520 not 387(2931) ; 387(2931)*
g3521 not 389(3021) ; 389(3021)*
g3522 not 390(2934) ; 390(2934)*
g3523 not 392(3022) ; 392(3022)*
g3524 not 393(2937) ; 393(2937)*
g3525 not 395(3023) ; 395(3023)*
g3526 not 396(2941) ; 396(2941)*
g3527 not 293(3285) ; 293(3285)*
g3528 not 294(3223) ; 294(3223)*
g3529 not 322(3302) ; 322(3302)*
g3530 not 323(3238) ; 323(3238)*
g3531 not 308(3346) ; 308(3346)*
g3532 not 309(3275) ; 309(3275)*
g3533 not 311(3349) ; 311(3349)*
g3534 not 312(3279) ; 312(3279)*
g3535 not 314(3350) ; 314(3350)*
g3536 not 315(3281) ; 315(3281)*
g3537 not 317(3351) ; 317(3351)*
g3538 not 318(3283) ; 318(3283)*
g3539 not 325(3358) ; 325(3358)*
g3540 not 326(3294) ; 326(3294)*
g3541 not 328(3361) ; 328(3361)*
g3542 not 329(3298) ; 329(3298)*
g3543 not 331(3364) ; 331(3364)*
g3544 not 332(3304) ; 332(3304)*
g3545 not 334(3362) ; 334(3362)*
g3546 not 335(3300) ; 335(3300)*
g3547 not 342(3330) ; 342(3330)*
g3548 not 343(3258) ; 343(3258)*
g3549 not 357(3376) ; 357(3376)*
g3550 not 358(3320) ; 358(3320)*
g3551 not 360(3379) ; 360(3379)*
g3552 not 361(3324) ; 361(3324)*
g3553 not 363(3380) ; 363(3380)*
g3554 not 364(3326) ; 364(3326)*
g3555 not 366(3381) ; 366(3381)*
g3556 not 367(3328) ; 367(3328)*
g3557 not 4528(206) ; 4528(206)*
g3558 not 1496(173) ; 1496(173)*
g3559 not 12(3) ; 12(3)*
g3560 not 9(2) ; 9(2)*
g3561 not 2207(272) ; 2207(272)*
g3562 not 1198(299) ; 1198(299)*
g3563 not 1519(374) ; 1519(374)*
g3564 not 6511(429) ; 6511(429)*
g3565 not 6518(558) ; 6518(558)*
g3566 not 5175(372) ; 5175(372)*
g3567 not 5182(563) ; 5182(563)*
g3568 not 4873(373) ; 4873(373)*
g3569 not 4880(566) ; 4880(566)*
g3570 not 4913(497) ; 4913(497)*
g3571 not 4920(565) ; 4920(565)*
g3572 not 5183(498) ; 5183(498)*
g3573 not 5190(562) ; 5190(562)*
g3574 not 5178(399) ; 5178(399)*
g3575 not 5181(494) ; 5181(494)*
g3576 not 4876(401) ; 4876(401)*
g3577 not 4879(495) ; 4879(495)*
g3578 not 1005(721) ; 1005(721)*
g3579 not 1006(602) ; 1006(602)*
g3580 not 763(723) ; 763(723)*
g3581 not 764(603) ; 764(603)*
g3582 not 6551(599) ; 6551(599)*
g3583 not 6558(556) ; 6558(556)*
g3584 not 6514(397) ; 6514(397)*
g3585 not 6517(598) ; 6517(598)*
g3586 not 5186(398) ; 5186(398)*
g3587 not 5189(607) ; 5189(607)*
g3588 not 4916(400) ; 4916(400)*
g3589 not 4919(605) ; 4919(605)*
g3590 not 3168(828) ; 3168(828)*
g3591 not 3169(597) ; 3169(597)*
g3592 not 737(854) ; 737(854)*
g3593 not 2241(257) ; 2241(257)*
g3594 not 2213(268) ; 2213(268)*
g3595 not 1399(820) ; 1399(820)*
g3596 not 885(832) ; 885(832)*
g3597 not 886(604) ; 886(604)*
g3598 not 1017(831) ; 1017(831)*
g3599 not 1018(606) ; 1018(606)*
g3600 not 1464(285) ; 1464(285)*
g3601 not 2933(861) ; 2933(861)*
g3602 not 6554(396) ; 6554(396)*
g3603 not 6557(741) ; 6557(741)*
g3604 not 4422(215) ; 4422(215)*
g3605 not 3821(1034) ; 3821(1034)*
g3606 not 4396(225) ; 4396(225)*
g3607 not 2179(977) ; 2179(977)*
g3608 not 3731(235) ; 3731(235)*
g3609 not 2091(969) ; 2091(969)*
g3610 not 5396(1084) ; 5396(1084)*
g3611 not 5399(466) ; 5399(466)*
g3612 not 5748(1085) ; 5748(1085)*
g3613 not 5751(467) ; 5751(467)*
g3614 not 5756(1086) ; 5756(1086)*
g3615 not 5759(469) ; 5759(469)*
g3616 not 5404(1087) ; 5404(1087)*
g3617 not 5407(470) ; 5407(470)*
g3618 not 5412(1076) ; 5412(1076)*
g3619 not 5415(472) ; 5415(472)*
g3620 not 5764(1075) ; 5764(1075)*
g3621 not 5767(473) ; 5767(473)*
g3622 not 5772(1078) ; 5772(1078)*
g3623 not 5775(474) ; 5775(474)*
g3624 not 5452(1077) ; 5452(1077)*
g3625 not 5455(475) ; 5455(475)*
g3626 not 5420(1082) ; 5420(1082)*
g3627 not 5423(478) ; 5423(478)*
g3628 not 5780(1081) ; 5780(1081)*
g3629 not 5783(479) ; 5783(479)*
g3630 not 5788(964) ; 5788(964)*
g3631 not 5791(480) ; 5791(480)*
g3632 not 5428(963) ; 5428(963)*
g3633 not 5431(481) ; 5431(481)*
g3634 not 5436(961) ; 5436(961)*
g3635 not 5439(484) ; 5439(484)*
g3636 not 5796(960) ; 5796(960)*
g3637 not 5799(485) ; 5799(485)*
g3638 not 5804(958) ; 5804(958)*
g3639 not 5807(486) ; 5807(486)*
g3640 not 5444(957) ; 5444(957)*
g3641 not 5447(487) ; 5447(487)*
g3642 not 5460(967) ; 5460(967)*
g3643 not 5463(489) ; 5463(489)*
g3644 not 7463(913) ; 7463(913)*
g3645 not 7470(915) ; 7470(915)*
g3646 not 5812(966) ; 5812(966)*
g3647 not 5815(491) ; 5815(491)*
g3648 not 6711(772) ; 6711(772)*
g3649 not 6718(921) ; 6718(921)*
g3650 not 777(370) ; 777(370)*
g3651 not 915(1029) ; 915(1029)*
g3652 not 6714(775) ; 6714(775)*
g3653 not 6717(916) ; 6717(916)*
g3654 not 4884(1105) ; 4884(1105)*
g3655 not 4887(500) ; 4887(500)*
g3656 not 5194(1106) ; 5194(1106)*
g3657 not 5197(501) ; 5197(501)*
g3658 not 5202(1089) ; 5202(1089)*
g3659 not 5205(502) ; 5205(502)*
g3660 not 4892(1090) ; 4892(1090)*
g3661 not 4895(503) ; 4895(503)*
g3662 not 5218(1095) ; 5218(1095)*
g3663 not 5221(505) ; 5221(505)*
g3664 not 4908(1096) ; 4908(1096)*
g3665 not 4911(507) ; 4911(507)*
g3666 not 4924(1099) ; 4924(1099)*
g3667 not 4927(508) ; 4927(508)*
g3668 not 6687(943) ; 6687(943)*
g3669 not 6694(945) ; 6694(945)*
g3670 not 5226(1100) ; 5226(1100)*
g3671 not 5229(510) ; 5229(510)*
g3672 not 7293(953) ; 7293(953)*
g3673 not 7300(946) ; 7300(946)*
g3674 not 5315(965) ; 5315(965)*
g3675 not 5322(955) ; 5322(955)*
g3676 not 4900(1093) ; 4900(1093)*
g3677 not 4903(671) ; 4903(671)*
g3678 not 5210(1094) ; 5210(1094)*
g3679 not 5213(672) ; 5213(672)*
g3680 not 7249(1024) ; 7249(1024)*
g3681 not 7256(1022) ; 7256(1022)*
g3682 not 3210(1026) ; 3210(1026)*
g3683 not 3211(827) ; 3211(827)*
g3684 not 5242(917) ; 5242(917)*
g3685 not 5245(830) ; 5245(830)*
g3686 not 5234(918) ; 5234(918)*
g3687 not 5237(720) ; 5237(720)*
g3688 not 5305(845) ; 5305(845)*
g3689 not 5312(1061) ; 5312(1061)*
g3690 not 5308(846) ; 5308(846)*
g3691 not 5311(1060) ; 5311(1060)*
g3692 not 5271(863) ; 5271(863)*
g3693 not 5278(1103) ; 5278(1103)*
g3694 not 5274(864) ; 5274(864)*
g3695 not 5277(1102) ; 5277(1102)*
g3696 not 6856(1327) ; 6856(1327)*
g3697 not 6859(431) ; 6859(431)*
g3698 not 6570(1329) ; 6570(1329)*
g3699 not 6573(432) ; 6573(432)*
g3700 not 6578(1350) ; 6578(1350)*
g3701 not 6581(433) ; 6581(433)*
g3702 not 6864(1352) ; 6864(1352)*
g3703 not 6867(434) ; 6867(434)*
g3704 not 6586(1378) ; 6586(1378)*
g3705 not 6589(435) ; 6589(435)*
g3706 not 6872(1377) ; 6872(1377)*
g3707 not 6875(436) ; 6875(436)*
g3708 not 6912(1374) ; 6912(1374)*
g3709 not 6915(437) ; 6915(437)*
g3710 not 6594(1375) ; 6594(1375)*
g3711 not 6597(438) ; 6597(438)*
g3712 not 6880(1361) ; 6880(1361)*
g3713 not 6883(439) ; 6883(439)*
g3714 not 6602(1359) ; 6602(1359)*
g3715 not 6605(440) ; 6605(440)*
g3716 not 6610(1266) ; 6610(1266)*
g3717 not 6613(441) ; 6613(441)*
g3718 not 6888(1267) ; 6888(1267)*
g3719 not 6891(442) ; 6891(442)*
g3720 not 6896(1302) ; 6896(1302)*
g3721 not 6899(443) ; 6899(443)*
g3722 not 6618(1303) ; 6618(1303)*
g3723 not 6621(444) ; 6621(444)*
g3724 not 6904(1296) ; 6904(1296)*
g3725 not 6907(445) ; 6907(445)*
g3726 not 6626(1297) ; 6626(1297)*
g3727 not 6629(446) ; 6629(446)*
g3728 not 6634(1275) ; 6634(1275)*
g3729 not 6637(447) ; 6637(447)*
g3730 not 6920(1276) ; 6920(1276)*
g3731 not 6923(448) ; 6923(448)*
g3732 not 5988(1290) ; 5988(1290)*
g3733 not 5991(449) ; 5991(449)*
g3734 not 5868(1291) ; 5868(1291)*
g3735 not 5871(450) ; 5871(450)*
g3736 not 5876(1259) ; 5876(1259)*
g3737 not 5879(451) ; 5879(451)*
g3738 not 5996(1260) ; 5996(1260)*
g3739 not 5999(452) ; 5999(452)*
g3740 not 6004(1254) ; 6004(1254)*
g3741 not 6007(453) ; 6007(453)*
g3742 not 5884(1255) ; 5884(1255)*
g3743 not 5887(454) ; 5887(454)*
g3744 not 6044(1251) ; 6044(1251)*
g3745 not 6047(455) ; 6047(455)*
g3746 not 5892(1250) ; 5892(1250)*
g3747 not 5895(456) ; 5895(456)*
g3748 not 5900(1288) ; 5900(1288)*
g3749 not 5903(457) ; 5903(457)*
g3750 not 6012(1287) ; 6012(1287)*
g3751 not 6015(458) ; 6015(458)*
g3752 not 6020(1395) ; 6020(1395)*
g3753 not 6023(459) ; 6023(459)*
g3754 not 5908(1394) ; 5908(1394)*
g3755 not 5911(460) ; 5911(460)*
g3756 not 5916(1390) ; 5916(1390)*
g3757 not 5919(461) ; 5919(461)*
g3758 not 6028(1389) ; 6028(1389)*
g3759 not 6031(462) ; 6031(462)*
g3760 not 6036(1383) ; 6036(1383)*
g3761 not 6039(463) ; 6039(463)*
g3762 not 5924(1382) ; 5924(1382)*
g3763 not 5927(464) ; 5927(464)*
g3764 not 7497(868) ; 7497(868)*
g3765 not 7504(1150) ; 7504(1150)*
g3766 not 6367(869) ; 6367(869)*
g3767 not 6374(1420) ; 6374(1420)*
g3768 not 5393(352) ; 5393(352)*
g3769 not 5400(1439) ; 5400(1439)*
g3770 not 5745(353) ; 5745(353)*
g3771 not 5752(1440) ; 5752(1440)*
g3772 not 7500(873) ; 7500(873)*
g3773 not 7503(1146) ; 7503(1146)*
g3774 not 6375(874) ; 6375(874)*
g3775 not 6382(1421) ; 6382(1421)*
g3776 not 5753(354) ; 5753(354)*
g3777 not 5760(1441) ; 5760(1441)*
g3778 not 5401(355) ; 5401(355)*
g3779 not 5408(1442) ; 5408(1442)*
g3780 not 6383(880) ; 6383(880)*
g3781 not 6390(1424) ; 6390(1424)*
g3782 not 7487(881) ; 7487(881)*
g3783 not 7494(1164) ; 7494(1164)*
g3784 not 5409(356) ; 5409(356)*
g3785 not 5416(1431) ; 5416(1431)*
g3786 not 5761(357) ; 5761(357)*
g3787 not 5768(1430) ; 5768(1430)*
g3788 not 5769(358) ; 5769(358)*
g3789 not 5776(1433) ; 5776(1433)*
g3790 not 5449(359) ; 5449(359)*
g3791 not 5456(1432) ; 5456(1432)*
g3792 not 7490(887) ; 7490(887)*
g3793 not 7493(1155) ; 7493(1155)*
g3794 not 6423(888) ; 6423(888)*
g3795 not 6430(1425) ; 6430(1425)*
g3796 not 7479(890) ; 7479(890)*
g3797 not 7486(1173) ; 7486(1173)*
g3798 not 6391(891) ; 6391(891)*
g3799 not 6398(1428) ; 6398(1428)*
g3800 not 5417(360) ; 5417(360)*
g3801 not 5424(1437) ; 5424(1437)*
g3802 not 5777(361) ; 5777(361)*
g3803 not 5784(1436) ; 5784(1436)*
g3804 not 5785(362) ; 5785(362)*
g3805 not 5792(1243) ; 5792(1243)*
g3806 not 5425(363) ; 5425(363)*
g3807 not 5432(1242) ; 5432(1242)*
g3808 not 6399(897) ; 6399(897)*
g3809 not 6406(1230) ; 6406(1230)*
g3810 not 7482(898) ; 7482(898)*
g3811 not 7485(1166) ; 7485(1166)*
g3812 not 7471(902) ; 7471(902)*
g3813 not 7478(1181) ; 7478(1181)*
g3814 not 6407(903) ; 6407(903)*
g3815 not 6414(1229) ; 6414(1229)*
g3816 not 5433(364) ; 5433(364)*
g3817 not 5440(1240) ; 5440(1240)*
g3818 not 5793(365) ; 5793(365)*
g3819 not 5800(1239) ; 5800(1239)*
g3820 not 5801(366) ; 5801(366)*
g3821 not 5808(1237) ; 5808(1237)*
g3822 not 5441(367) ; 5441(367)*
g3823 not 5448(1236) ; 5448(1236)*
g3824 not 6415(907) ; 6415(907)*
g3825 not 6422(1226) ; 6422(1226)*
g3826 not 7474(908) ; 7474(908)*
g3827 not 7477(1174) ; 7477(1174)*
g3828 not 5457(368) ; 5457(368)*
g3829 not 5464(1246) ; 5464(1246)*
g3830 not 6431(914) ; 6431(914)*
g3831 not 6438(1233) ; 6438(1233)*
g3832 not 5809(369) ; 5809(369)*
g3833 not 5816(1245) ; 5816(1245)*
g3834 not 7466(771) ; 7466(771)*
g3835 not 7469(1186) ; 7469(1186)*
g3836 not 6719(1202) ; 6719(1202)*
g3837 not 6720(1189) ; 6720(1189)*
g3838 not 6703(927) ; 6703(927)*
g3839 not 6710(1213) ; 6710(1213)*
g3840 not 6519(928) ; 6519(928)*
g3841 not 6526(1418) ; 6526(1418)*
g3842 not 4881(375) ; 4881(375)*
g3843 not 4888(1460) ; 4888(1460)*
g3844 not 5191(376) ; 5191(376)*
g3845 not 5198(1461) ; 5198(1461)*
g3846 not 5199(377) ; 5199(377)*
g3847 not 5206(1444) ; 5206(1444)*
g3848 not 4889(378) ; 4889(378)*
g3849 not 4896(1445) ; 4896(1445)*
g3850 not 6527(932) ; 6527(932)*
g3851 not 6534(1408) ; 6534(1408)*
g3852 not 6706(933) ; 6706(933)*
g3853 not 6709(1206) ; 6709(1206)*
g3854 not 5215(379) ; 5215(379)*
g3855 not 5222(1450) ; 5222(1450)*
g3856 not 6543(937) ; 6543(937)*
g3857 not 6550(1412) ; 6550(1412)*
g3858 not 6698(938) ; 6698(938)*
g3859 not 6701(1281) ; 6701(1281)*
g3860 not 4905(380) ; 4905(380)*
g3861 not 4912(1451) ; 4912(1451)*
g3862 not 4921(381) ; 4921(381)*
g3863 not 4928(1454) ; 4928(1454)*
g3864 not 6559(944) ; 6559(944)*
g3865 not 6566(1414) ; 6566(1414)*
g3866 not 5223(382) ; 5223(382)*
g3867 not 5230(1455) ; 5230(1455)*
g3868 not 6690(780) ; 6690(780)*
g3869 not 6693(1222) ; 6693(1222)*
g3870 not 7296(811) ; 7296(811)*
g3871 not 7299(1232) ; 7299(1232)*
g3872 not 6418(947) ; 6418(947)*
g3873 not 6421(1180) ; 6421(1180)*
g3874 not 7304(948) ; 7304(948)*
g3875 not 7307(1228) ; 7307(1228)*
g3876 not 7301(949) ; 7301(949)*
g3877 not 7308(1227) ; 7308(1227)*
g3878 not 6410(950) ; 6410(950)*
g3879 not 6413(1175) ; 6413(1175)*
g3880 not 6402(951) ; 6402(951)*
g3881 not 6405(1172) ; 6405(1172)*
g3882 not 7312(952) ; 7312(952)*
g3883 not 7315(1427) ; 7315(1427)*
g3884 not 6434(954) ; 6434(954)*
g3885 not 6437(1187) ; 6437(1187)*
g3886 not 5318(816) ; 5318(816)*
g3887 not 5321(1244) ; 5321(1244)*
g3888 not 5326(956) ; 5326(956)*
g3889 not 5329(1238) ; 5329(1238)*
g3890 not 5323(959) ; 5323(959)*
g3891 not 5330(1235) ; 5330(1235)*
g3892 not 5334(962) ; 5334(962)*
g3893 not 5337(1435) ; 5337(1435)*
g3894 not 7224(1270) ; 7224(1270)*
g3895 not 7227(1358) ; 7227(1358)*
g3896 not 7205(1273) ; 7205(1273)*
g3897 not 7212(1277) ; 7212(1277)*
g3898 not 6721(1274) ; 6721(1274)*
g3899 not 6728(1278) ; 6728(1278)*
g3900 not 4897(548) ; 4897(548)*
g3901 not 4904(1448) ; 4904(1448)*
g3902 not 5207(549) ; 5207(549)*
g3903 not 5214(1449) ; 5214(1449)*
g3904 not 6695(983) ; 6695(983)*
g3905 not 6702(1216) ; 6702(1216)*
g3906 not 6535(984) ; 6535(984)*
g3907 not 6542(1410) ; 6542(1410)*
g3908 not 7265(1285) ; 7265(1285)*
g3909 not 7272(1399) ; 7272(1399)*
g3910 not 6463(1309) ; 6463(1309)*
g3911 not 6470(1357) ; 6470(1357)*
g3912 not 6495(1311) ; 6495(1311)*
g3913 not 6502(1371) ; 6502(1371)*
g3914 not 7551(1316) ; 7551(1316)*
g3915 not 7558(1341) ; 7558(1341)*
g3916 not 7401(1318) ; 7401(1318)*
g3917 not 7408(1391) ; 7408(1391)*
g3918 not 7393(1319) ; 7393(1319)*
g3919 not 7400(1398) ; 7400(1398)*
g3920 not 7409(1321) ; 7409(1321)*
g3921 not 7416(1386) ; 7416(1386)*
g3922 not 7507(1002) ; 7507(1002)*
g3923 not 7514(1326) ; 7514(1326)*
g3924 not 7510(1003) ; 7510(1003)*
g3925 not 7513(1325) ; 7513(1325)*
g3926 not 7239(1005) ; 7239(1005)*
g3927 not 7246(1355) ; 7246(1355)*
g3928 not 6439(1333) ; 6439(1333)*
g3929 not 6446(1332) ; 6446(1332)*
g3930 not 6447(1335) ; 6447(1335)*
g3931 not 6454(1354) ; 6454(1354)*
g3932 not 6455(1337) ; 6455(1337)*
g3933 not 6462(1380) ; 6462(1380)*
g3934 not 7242(1018) ; 7242(1018)*
g3935 not 7245(1331) ; 7245(1331)*
g3936 not 7252(825) ; 7252(825)*
g3937 not 7255(1364) ; 7255(1364)*
g3938 not 6765(1365) ; 6765(1365)*
g3939 not 6772(1363) ; 6772(1363)*
g3940 not 5239(719) ; 5239(719)*
g3941 not 5246(1194) ; 5246(1194)*
g3942 not 5231(561) ; 5231(561)*
g3943 not 5238(1195) ; 5238(1195)*
g3944 not 7232(1033) ; 7232(1033)*
g3945 not 7235(1381) ; 7235(1381)*
g3946 not 7229(1037) ; 7229(1037)*
g3947 not 7236(1372) ; 7236(1372)*
g3948 not 7260(1040) ; 7260(1040)*
g3949 not 7263(1393) ; 7263(1393)*
g3950 not 7257(1043) ; 7257(1043)*
g3951 not 7264(1387) ; 7264(1387)*
g3952 not 7428(1404) ; 7428(1404)*
g3953 not 7431(1401) ; 7431(1401)*
g3954 not 3682(839) ; 3682(839)*
g3955 not 4389(1405) ; 4389(1405)*
g3956 not 5284(1051) ; 5284(1051)*
g3957 not 5287(1413) ; 5287(1413)*
g3958 not 5300(1052) ; 5300(1052)*
g3959 not 5303(1417) ; 5303(1417)*
g3960 not 6530(1053) ; 6530(1053)*
g3961 not 6533(1212) ; 6533(1212)*
g3962 not 5289(1054) ; 5289(1054)*
g3963 not 5296(1411) ; 5296(1411)*
g3964 not 6538(1055) ; 6538(1055)*
g3965 not 6541(1282) ; 6541(1282)*
g3966 not 5292(1056) ; 5292(1056)*
g3967 not 5295(1409) ; 5295(1409)*
g3968 not 6546(1057) ; 6546(1057)*
g3969 not 6549(1215) ; 6549(1215)*
g3970 not 5281(1058) ; 5281(1058)*
g3971 not 5288(1406) ; 5288(1406)*
g3972 not 6562(1059) ; 6562(1059)*
g3973 not 6565(1223) ; 6565(1223)*
g3974 not 5313(1416) ; 5313(1416)*
g3975 not 5314(1415) ; 5314(1415)*
g3976 not 5297(1062) ; 5297(1062)*
g3977 not 5304(1407) ; 5304(1407)*
g3978 not 6522(1063) ; 6522(1063)*
g3979 not 6525(1207) ; 6525(1207)*
g3980 not 7327(1064) ; 7327(1064)*
g3981 not 7334(1422) ; 7334(1422)*
g3982 not 6370(1065) ; 6370(1065)*
g3983 not 6373(1147) ; 6373(1147)*
g3984 not 6378(1066) ; 6378(1066)*
g3985 not 6381(1151) ; 6381(1151)*
g3986 not 7330(1067) ; 7330(1067)*
g3987 not 7333(1419) ; 7333(1419)*
g3988 not 7317(1068) ; 7317(1068)*
g3989 not 7324(1426) ; 7324(1426)*
g3990 not 6386(1069) ; 6386(1069)*
g3991 not 6389(1154) ; 6389(1154)*
g3992 not 6426(1070) ; 6426(1070)*
g3993 not 6429(1165) ; 6429(1165)*
g3994 not 7320(1071) ; 7320(1071)*
g3995 not 7323(1423) ; 7323(1423)*
g3996 not 7309(1072) ; 7309(1072)*
g3997 not 7316(1231) ; 7316(1231)*
g3998 not 6394(1073) ; 6394(1073)*
g3999 not 6397(1167) ; 6397(1167)*
g4000 not 5339(1074) ; 5339(1074)*
g4001 not 5346(1434) ; 5346(1434)*
g4002 not 5342(1079) ; 5342(1079)*
g4003 not 5345(1429) ; 5345(1429)*
g4004 not 5331(1080) ; 5331(1080)*
g4005 not 5338(1241) ; 5338(1241)*
g4006 not 5349(1083) ; 5349(1083)*
g4007 not 5356(1443) ; 5356(1443)*
g4008 not 5352(1088) ; 5352(1088)*
g4009 not 5355(1438) ; 5355(1438)*
g4010 not 5266(1091) ; 5266(1091)*
g4011 not 5269(1459) ; 5269(1459)*
g4012 not 5255(1092) ; 5255(1092)*
g4013 not 5262(1452) ; 5262(1452)*
g4014 not 5258(1097) ; 5258(1097)*
g4015 not 5261(1447) ; 5261(1447)*
g4016 not 5247(1098) ; 5247(1098)*
g4017 not 5254(1456) ; 5254(1456)*
g4018 not 5250(1101) ; 5250(1101)*
g4019 not 5253(1453) ; 5253(1453)*
g4020 not 5279(1458) ; 5279(1458)*
g4021 not 5280(1457) ; 5280(1457)*
g4022 not 5263(1104) ; 5263(1104)*
g4023 not 5270(1446) ; 5270(1446)*
g4024 not 6853(318) ; 6853(318)*
g4025 not 6860(1665) ; 6860(1665)*
g4026 not 6567(319) ; 6567(319)*
g4027 not 6574(1667) ; 6574(1667)*
g4028 not 6575(320) ; 6575(320)*
g4029 not 6582(1688) ; 6582(1688)*
g4030 not 6861(321) ; 6861(321)*
g4031 not 6868(1690) ; 6868(1690)*
g4032 not 6583(322) ; 6583(322)*
g4033 not 6590(1707) ; 6590(1707)*
g4034 not 6869(323) ; 6869(323)*
g4035 not 6876(1706) ; 6876(1706)*
g4036 not 6909(324) ; 6909(324)*
g4037 not 6916(1703) ; 6916(1703)*
g4038 not 6591(325) ; 6591(325)*
g4039 not 6598(1704) ; 6598(1704)*
g4040 not 6877(326) ; 6877(326)*
g4041 not 6884(1694) ; 6884(1694)*
g4042 not 6599(327) ; 6599(327)*
g4043 not 6606(1692) ; 6606(1692)*
g4044 not 6607(328) ; 6607(328)*
g4045 not 6614(1602) ; 6614(1602)*
g4046 not 6885(329) ; 6885(329)*
g4047 not 6892(1603) ; 6892(1603)*
g4048 not 6893(330) ; 6893(330)*
g4049 not 6900(1635) ; 6900(1635)*
g4050 not 6615(331) ; 6615(331)*
g4051 not 6622(1636) ; 6622(1636)*
g4052 not 6901(332) ; 6901(332)*
g4053 not 6908(1630) ; 6908(1630)*
g4054 not 6623(333) ; 6623(333)*
g4055 not 6630(1631) ; 6630(1631)*
g4056 not 6631(334) ; 6631(334)*
g4057 not 6638(1612) ; 6638(1612)*
g4058 not 6917(335) ; 6917(335)*
g4059 not 6924(1613) ; 6924(1613)*
g4060 not 5985(336) ; 5985(336)*
g4061 not 5992(1625) ; 5992(1625)*
g4062 not 5865(337) ; 5865(337)*
g4063 not 5872(1626) ; 5872(1626)*
g4064 not 5873(338) ; 5873(338)*
g4065 not 5880(1596) ; 5880(1596)*
g4066 not 5993(339) ; 5993(339)*
g4067 not 6000(1597) ; 6000(1597)*
g4068 not 6001(340) ; 6001(340)*
g4069 not 6008(1592) ; 6008(1592)*
g4070 not 5881(341) ; 5881(341)*
g4071 not 5888(1593) ; 5888(1593)*
g4072 not 6041(342) ; 6041(342)*
g4073 not 6048(1589) ; 6048(1589)*
g4074 not 5889(343) ; 5889(343)*
g4075 not 5896(1588) ; 5896(1588)*
g4076 not 5897(344) ; 5897(344)*
g4077 not 5904(1623) ; 5904(1623)*
g4078 not 6009(345) ; 6009(345)*
g4079 not 6016(1622) ; 6016(1622)*
g4080 not 6017(346) ; 6017(346)*
g4081 not 6024(1718) ; 6024(1718)*
g4082 not 5905(347) ; 5905(347)*
g4083 not 5912(1717) ; 5912(1717)*
g4084 not 5913(348) ; 5913(348)*
g4085 not 5920(1715) ; 5920(1715)*
g4086 not 6025(349) ; 6025(349)*
g4087 not 6032(1714) ; 6032(1714)*
g4088 not 6033(350) ; 6033(350)*
g4089 not 6040(1710) ; 6040(1710)*
g4090 not 5921(351) ; 5921(351)*
g4091 not 5928(1709) ; 5928(1709)*
g4092 not 7505(1511) ; 7505(1511)*
g4093 not 7506(1507) ; 7506(1507)*
g4094 not 2954(1740) ; 2954(1740)*
g4095 not 2955(1508) ; 2955(1508)*
g4096 not 1544(1148) ; 1544(1148)*
g4097 not 1545(1509) ; 1545(1509)*
g4098 not 1793(1149) ; 1793(1149)*
g4099 not 1794(1510) ; 1794(1510)*
g4100 not 2963(1741) ; 2963(1741)*
g4101 not 2964(1512) ; 2964(1512)*
g4102 not 1803(1152) ; 1803(1152)*
g4103 not 1804(1513) ; 1804(1513)*
g4104 not 1554(1153) ; 1554(1153)*
g4105 not 1555(1514) ; 1555(1514)*
g4106 not 2971(1744) ; 2971(1744)*
g4107 not 2972(1515) ; 2972(1515)*
g4108 not 7495(1523) ; 7495(1523)*
g4109 not 7496(1516) ; 7496(1516)*
g4110 not 1571(1156) ; 1571(1156)*
g4111 not 1572(1517) ; 1572(1517)*
g4112 not 1820(1157) ; 1820(1157)*
g4113 not 1821(1518) ; 1821(1518)*
g4114 not 1848(1160) ; 1848(1160)*
g4115 not 1849(1521) ; 1849(1521)*
g4116 not 1685(1163) ; 1685(1163)*
g4117 not 1686(1522) ; 1686(1522)*
g4118 not 3016(1745) ; 3016(1745)*
g4119 not 3017(1524) ; 3017(1524)*
g4120 not 4547(1532) ; 4547(1532)*
g4121 not 4548(1525) ; 4548(1525)*
g4122 not 2980(1748) ; 2980(1748)*
g4123 not 2981(1526) ; 2981(1526)*
g4124 not 1596(1168) ; 1596(1168)*
g4125 not 1597(1527) ; 1597(1527)*
g4126 not 1857(1169) ; 1857(1169)*
g4127 not 1858(1528) ; 1858(1528)*
g4128 not 1867(1170) ; 1867(1170)*
g4129 not 1868(1529) ; 1868(1529)*
g4130 not 1607(1171) ; 1607(1171)*
g4131 not 1608(1530) ; 1608(1530)*
g4132 not 2990(1579) ; 2990(1579)*
g4133 not 2991(1531) ; 2991(1531)*
g4134 not 4538(1540) ; 4538(1540)*
g4135 not 4539(1533) ; 4539(1533)*
g4136 not 2999(1578) ; 2999(1578)*
g4137 not 3000(1534) ; 3000(1534)*
g4138 not 1628(1176) ; 1628(1176)*
g4139 not 1629(1535) ; 1629(1535)*
g4140 not 1883(1177) ; 1883(1177)*
g4141 not 1884(1536) ; 1884(1536)*
g4142 not 1901(1178) ; 1901(1178)*
g4143 not 1902(1537) ; 1902(1537)*
g4144 not 1653(1179) ; 1653(1179)*
g4145 not 1654(1538) ; 1654(1538)*
g4146 not 3007(1575) ; 3007(1575)*
g4147 not 3008(1539) ; 3008(1539)*
g4148 not 1693(1184) ; 1693(1184)*
g4149 not 1694(1542) ; 1694(1542)*
g4150 not 4529(1545) ; 4529(1545)*
g4151 not 4530(1185) ; 4530(1185)*
g4152 not 3019(1581) ; 3019(1581)*
g4153 not 3020(1543) ; 3020(1543)*
g4154 not 1919(1188) ; 1919(1188)*
g4155 not 1920(1544) ; 1920(1544)*
g4156 not 912(1550) ; 912(1550)*
g4157 not 906(1554) ; 906(1554)*
g4158 not 1121(1552) ; 1121(1552)*
g4159 not 1112(1553) ; 1112(1553)*
g4160 not 3520(1564) ; 3520(1564)*
g4161 not 3521(1557) ; 3521(1557)*
g4162 not 3174(1738) ; 3174(1738)*
g4163 not 3175(1558) ; 3175(1558)*
g4164 not 790(1208) ; 790(1208)*
g4165 not 791(1559) ; 791(1559)*
g4166 not 1024(1209) ; 1024(1209)*
g4167 not 1025(1560) ; 1025(1560)*
g4168 not 1036(1210) ; 1036(1210)*
g4169 not 1037(1561) ; 1037(1561)*
g4170 not 803(1211) ; 803(1211)*
g4171 not 804(1562) ; 804(1562)*
g4172 not 3184(1729) ; 3184(1729)*
g4173 not 3185(1563) ; 3185(1563)*
g4174 not 1072(1214) ; 1072(1214)*
g4175 not 1073(1565) ; 1073(1565)*
g4176 not 3201(1733) ; 3201(1733)*
g4177 not 3202(1566) ; 3202(1566)*
g4178 not 3511(1567) ; 3511(1567)*
g4179 not 3512(1616) ; 3512(1616)*
g4180 not 851(1217) ; 851(1217)*
g4181 not 852(1568) ; 852(1568)*
g4182 not 893(1220) ; 893(1220)*
g4183 not 894(1570) ; 894(1570)*
g4184 not 3502(1573) ; 3502(1573)*
g4185 not 3503(1221) ; 3503(1221)*
g4186 not 3213(1735) ; 3213(1735)*
g4187 not 3214(1571) ; 3214(1571)*
g4188 not 1091(1224) ; 1091(1224)*
g4189 not 1092(1572) ; 1092(1572)*
g4190 not 4224(1574) ; 4224(1574)*
g4191 not 4225(1225) ; 4225(1225)*
g4192 not 4233(1576) ; 4233(1576)*
g4193 not 4234(1577) ; 4234(1577)*
g4194 not 4242(1580) ; 4242(1580)*
g4195 not 4243(1747) ; 4243(1747)*
g4196 not 1261(1582) ; 1261(1582)*
g4197 not 1262(1234) ; 1262(1234)*
g4198 not 1270(1583) ; 1270(1583)*
g4199 not 1271(1584) ; 1271(1584)*
g4200 not 1279(1585) ; 1279(1585)*
g4201 not 1280(1751) ; 1280(1751)*
g4202 not 7276(1247) ; 7276(1247)*
g4203 not 7279(1595) ; 7279(1595)*
g4204 not 7420(1249) ; 7420(1249)*
g4205 not 7423(1687) ; 7423(1687)*
g4206 not 6792(1252) ; 6792(1252)*
g4207 not 6795(1591) ; 6795(1591)*
g4208 not 6789(1253) ; 6789(1253)*
g4209 not 6796(1590) ; 6796(1590)*
g4210 not 7380(1257) ; 7380(1257)*
g4211 not 7383(1685) ; 7383(1685)*
g4212 not 7273(1258) ; 7273(1258)*
g4213 not 7280(1586) ; 7280(1586)*
g4214 not 6802(1261) ; 6802(1261)*
g4215 not 6805(1624) ; 6805(1624)*
g4216 not 7372(1263) ; 7372(1263)*
g4217 not 7375(1682) ; 7375(1682)*
g4218 not 7286(1264) ; 7286(1264)*
g4219 not 7289(1628) ; 7289(1628)*
g4220 not 6740(1265) ; 6740(1265)*
g4221 not 6743(1693) ; 6743(1693)*
g4222 not 6474(1269) ; 6474(1269)*
g4223 not 6477(1639) ; 6477(1639)*
g4224 not 6506(1272) ; 6506(1272)*
g4225 not 6509(1649) ; 6509(1649)*
g4226 not 7208(978) ; 7208(978)*
g4227 not 7211(1609) ; 7211(1609)*
g4228 not 6724(979) ; 6724(979)*
g4229 not 6727(1611) ; 6727(1611)*
g4230 not 825(1279) ; 825(1279)*
g4231 not 826(1614) ; 826(1614)*
g4232 not 1053(1280) ; 1053(1280)*
g4233 not 1054(1615) ; 1054(1615)*
g4234 not 3193(1731) ; 3193(1731)*
g4235 not 3194(1617) ; 3194(1617)*
g4236 not 7388(1283) ; 7388(1283)*
g4237 not 7391(1662) ; 7391(1662)*
g4238 not 6781(1286) ; 6781(1286)*
g4239 not 6788(1719) ; 6788(1719)*
g4240 not 6799(1289) ; 6799(1289)*
g4241 not 6806(1598) ; 6806(1598)*
g4242 not 7364(1292) ; 7364(1292)*
g4243 not 7367(1681) ; 7367(1681)*
g4244 not 7283(1294) ; 7283(1294)*
g4245 not 7290(1600) ; 7290(1600)*
g4246 not 6732(1295) ; 6732(1295)*
g4247 not 6735(1634) ; 6735(1634)*
g4248 not 6490(1299) ; 6490(1299)*
g4249 not 6493(1647) ; 6493(1647)*
g4250 not 7216(1300) ; 7216(1300)*
g4251 not 7219(1638) ; 7219(1638)*
g4252 not 6729(1301) ; 6729(1301)*
g4253 not 6736(1629) ; 6736(1629)*
g4254 not 6482(1304) ; 6482(1304)*
g4255 not 6485(1678) ; 6485(1678)*
g4256 not 7213(1306) ; 7213(1306)*
g4257 not 7220(1633) ; 7220(1633)*
g4258 not 6471(1307) ; 6471(1307)*
g4259 not 6478(1604) ; 6478(1604)*
g4260 not 7570(1308) ; 7570(1308)*
g4261 not 7573(1643) ; 7573(1643)*
g4262 not 7567(1310) ; 7567(1310)*
g4263 not 7574(1640) ; 7574(1640)*
g4264 not 7578(1312) ; 7578(1312)*
g4265 not 7581(1677) ; 7581(1677)*
g4266 not 6487(1313) ; 6487(1313)*
g4267 not 6494(1632) ; 6494(1632)*
g4268 not 7562(1314) ; 7562(1314)*
g4269 not 7565(1679) ; 7565(1679)*
g4270 not 6503(1315) ; 6503(1315)*
g4271 not 6510(1607) ; 6510(1607)*
g4272 not 7515(1317) ; 7515(1317)*
g4273 not 7522(1660) ; 7522(1660)*
g4274 not 7526(1320) ; 7526(1320)*
g4275 not 7529(1661) ; 7529(1661)*
g4276 not 7518(1322) ; 7518(1322)*
g4277 not 7521(1652) ; 7521(1652)*
g4278 not 7523(1323) ; 7523(1323)*
g4279 not 7530(1657) ; 7530(1657)*
g4280 not 7385(1324) ; 7385(1324)*
g4281 not 7392(1618) ; 7392(1618)*
g4282 not 4552(1664) ; 4552(1664)*
g4283 not 4553(1663) ; 4553(1663)*
g4284 not 6755(1328) ; 6755(1328)*
g4285 not 6762(1689) ; 6762(1689)*
g4286 not 7247(1691) ; 7247(1691)*
g4287 not 7248(1668) ; 7248(1668)*
g4288 not 6442(1006) ; 6442(1006)*
g4289 not 6445(1670) ; 6445(1670)*
g4290 not 7585(1334) ; 7585(1334)*
g4291 not 7592(1674) ; 7592(1674)*
g4292 not 7588(1336) ; 7588(1336)*
g4293 not 7591(1671) ; 7591(1671)*
g4294 not 7575(1338) ; 7575(1338)*
g4295 not 7582(1646) ; 7582(1646)*
g4296 not 6479(1339) ; 6479(1339)*
g4297 not 6486(1637) ; 6486(1637)*
g4298 not 7559(1340) ; 7559(1340)*
g4299 not 7566(1648) ; 7566(1648)*
g4300 not 7554(1011) ; 7554(1011)*
g4301 not 7557(1651) ; 7557(1651)*
g4302 not 7541(1342) ; 7541(1342)*
g4303 not 7548(1683) ; 7548(1683)*
g4304 not 7361(1343) ; 7361(1343)*
g4305 not 7368(1627) ; 7368(1627)*
g4306 not 7369(1344) ; 7369(1344)*
g4307 not 7376(1599) ; 7376(1599)*
g4308 not 7544(1345) ; 7544(1345)*
g4309 not 7547(1680) ; 7547(1680)*
g4310 not 7531(1346) ; 7531(1346)*
g4311 not 7538(1686) ; 7538(1686)*
g4312 not 7377(1347) ; 7377(1347)*
g4313 not 7384(1594) ; 7384(1594)*
g4314 not 7534(1348) ; 7534(1348)*
g4315 not 7537(1684) ; 7537(1684)*
g4316 not 7417(1349) ; 7417(1349)*
g4317 not 7424(1587) ; 7424(1587)*
g4318 not 6758(1351) ; 6758(1351)*
g4319 not 6761(1666) ; 6761(1666)*
g4320 not 6450(1017) ; 6450(1017)*
g4321 not 6453(1673) ; 6453(1673)*
g4322 not 6466(1019) ; 6466(1019)*
g4323 not 6469(1642) ; 6469(1642)*
g4324 not 7221(1020) ; 7221(1020)*
g4325 not 7228(1606) ; 7228(1606)*
g4326 not 6737(1360) ; 6737(1360)*
g4327 not 6744(1601) ; 6744(1601)*
g4328 not 4201(1695) ; 4201(1695)*
g4329 not 4202(1362) ; 4202(1362)*
g4330 not 6768(1023) ; 6768(1023)*
g4331 not 6771(1697) ; 6771(1697)*
g4332 not 4973(1548) ; 4973(1548)*
g4333 not 4976(829) ; 4976(829)*
g4334 not 1156(1368) ; 1156(1368)*
g4335 not 1157(1699) ; 1157(1699)*
g4336 not 1152(1369) ; 1152(1369)*
g4337 not 1153(1700) ; 1153(1700)*
g4338 not 4932(1547) ; 4932(1547)*
g4339 not 4935(722) ; 4935(722)*
g4340 not 6498(1032) ; 6498(1032)*
g4341 not 6501(1645) ; 6501(1645)*
g4342 not 7237(1701) ; 7237(1701)*
g4343 not 7238(1708) ; 7238(1708)*
g4344 not 6748(1373) ; 6748(1373)*
g4345 not 6751(1705) ; 6751(1705)*
g4346 not 6745(1376) ; 6745(1376)*
g4347 not 6752(1702) ; 6752(1702)*
g4348 not 6458(1036) ; 6458(1036)*
g4349 not 6461(1676) ; 6461(1676)*
g4350 not 6776(1384) ; 6776(1384)*
g4351 not 6779(1713) ; 6779(1713)*
g4352 not 7412(1039) ; 7412(1039)*
g4353 not 7415(1659) ; 7415(1659)*
g4354 not 4210(1712) ; 4210(1712)*
g4355 not 4211(1716) ; 4211(1716)*
g4356 not 6773(1388) ; 6773(1388)*
g4357 not 6780(1711) ; 6780(1711)*
g4358 not 7404(1042) ; 7404(1042)*
g4359 not 7407(1654) ; 7407(1654)*
g4360 not 6784(1396) ; 6784(1396)*
g4361 not 6787(1621) ; 6787(1621)*
g4362 not 7396(1045) ; 7396(1045)*
g4363 not 7399(1656) ; 7399(1656)*
g4364 not 7268(1046) ; 7268(1046)*
g4365 not 7271(1620) ; 7271(1620)*
g4366 not 7425(1047) ; 7425(1047)*
g4367 not 7432(1724) ; 7432(1724)*
g4368 not 5932(1726) ; 5932(1726)*
g4369 not 5935(1402) ; 5935(1402)*
g4370 not 6052(1725) ; 6052(1725)*
g4371 not 6055(1403) ; 6055(1403)*
g4372 not 1238(1727) ; 1238(1727)*
g4373 not 1239(1734) ; 1239(1734)*
g4374 not 1256(1728) ; 1256(1728)*
g4375 not 1257(1737) ; 1257(1737)*
g4376 not 1247(1732) ; 1247(1732)*
g4377 not 1248(1730) ; 1248(1730)*
g4378 not 7335(1742) ; 7335(1742)*
g4379 not 7336(1739) ; 7336(1739)*
g4380 not 7325(1746) ; 7325(1746)*
g4381 not 7326(1743) ; 7326(1743)*
g4382 not 5347(1750) ; 5347(1750)*
g4383 not 5348(1749) ; 5348(1749)*
g4384 not 5357(1753) ; 5357(1753)*
g4385 not 5358(1752) ; 5358(1752)*
g4386 not 1233(1754) ; 1233(1754)*
g4387 not 1234(1760) ; 1234(1760)*
g4388 not 1224(1756) ; 1224(1756)*
g4389 not 1225(1755) ; 1225(1755)*
g4390 not 1215(1758) ; 1215(1758)*
g4391 not 1216(1757) ; 1216(1757)*
g4392 not 3227(1925) ; 3227(1925)*
g4393 not 3220(1761) ; 3220(1761)*
g4394 not 3843(1463) ; 3843(1463)*
g4395 not 3844(1762) ; 3844(1762)*
g4396 not 3281(1464) ; 3281(1464)*
g4397 not 3282(1763) ; 3282(1763)*
g4398 not 3293(1465) ; 3293(1465)*
g4399 not 3294(1764) ; 3294(1764)*
g4400 not 3854(1466) ; 3854(1466)*
g4401 not 3855(1765) ; 3855(1765)*
g4402 not 3312(1467) ; 3312(1467)*
g4403 not 3313(1766) ; 3313(1766)*
g4404 not 3872(1468) ; 3872(1468)*
g4405 not 3873(1767) ; 3873(1767)*
g4406 not 3987(1472) ; 3987(1472)*
g4407 not 3988(1770) ; 3988(1770)*
g4408 not 3342(1473) ; 3342(1473)*
g4409 not 3343(1771) ; 3343(1771)*
g4410 not 3897(1475) ; 3897(1475)*
g4411 not 3898(1772) ; 3898(1772)*
g4412 not 3351(1476) ; 3351(1476)*
g4413 not 3352(1773) ; 3352(1773)*
g4414 not 3363(1477) ; 3363(1477)*
g4415 not 3364(1774) ; 3364(1774)*
g4416 not 3909(1478) ; 3909(1478)*
g4417 not 3910(1775) ; 3910(1775)*
g4418 not 3930(1479) ; 3930(1479)*
g4419 not 3931(1776) ; 3931(1776)*
g4420 not 3379(1480) ; 3379(1480)*
g4421 not 3380(1777) ; 3380(1777)*
g4422 not 3955(1481) ; 3955(1481)*
g4423 not 3956(1778) ; 3956(1778)*
g4424 not 3397(1482) ; 3397(1482)*
g4425 not 3398(1779) ; 3398(1779)*
g4426 not 3415(1484) ; 3415(1484)*
g4427 not 3416(1781) ; 3416(1781)*
g4428 not 3995(1486) ; 3995(1486)*
g4429 not 3996(1782) ; 3996(1782)*
g4430 not 2587(1487) ; 2587(1487)*
g4431 not 2588(1783) ; 2588(1783)*
g4432 not 2341(1488) ; 2341(1488)*
g4433 not 2342(1784) ; 2342(1784)*
g4434 not 2352(1489) ; 2352(1489)*
g4435 not 2353(1785) ; 2353(1785)*
g4436 not 2598(1490) ; 2598(1490)*
g4437 not 2599(1786) ; 2599(1786)*
g4438 not 2616(1491) ; 2616(1491)*
g4439 not 2617(1787) ; 2617(1787)*
g4440 not 2370(1492) ; 2370(1492)*
g4441 not 2371(1788) ; 2371(1788)*
g4442 not 2732(1496) ; 2732(1496)*
g4443 not 2733(1791) ; 2733(1791)*
g4444 not 2398(1497) ; 2398(1497)*
g4445 not 2399(1792) ; 2399(1792)*
g4446 not 2407(1499) ; 2407(1499)*
g4447 not 2408(1793) ; 2408(1793)*
g4448 not 2641(1500) ; 2641(1500)*
g4449 not 2642(1794) ; 2642(1794)*
g4450 not 2653(1501) ; 2653(1501)*
g4451 not 2654(1795) ; 2654(1795)*
g4452 not 2418(1502) ; 2418(1502)*
g4453 not 2419(1796) ; 2419(1796)*
g4454 not 2434(1503) ; 2434(1503)*
g4455 not 2435(1797) ; 2435(1797)*
g4456 not 2674(1504) ; 2674(1504)*
g4457 not 2675(1798) ; 2675(1798)*
g4458 not 2699(1505) ; 2699(1505)*
g4459 not 2700(1799) ; 2700(1799)*
g4460 not 2452(1506) ; 2452(1506)*
g4461 not 2453(1800) ; 2453(1800)*
g4462 not 7281(1860) ; 7281(1860)*
g4463 not 7282(1865) ; 7282(1865)*
g4464 not 4350(1861) ; 4350(1861)*
g4465 not 4351(1917) ; 4351(1917)*
g4466 not 6797(1862) ; 6797(1862)*
g4467 not 6798(1863) ; 6798(1863)*
g4468 not 4306(1864) ; 4306(1864)*
g4469 not 4307(1915) ; 4307(1915)*
g4470 not 6807(1866) ; 6807(1866)*
g4471 not 6808(1879) ; 6808(1879)*
g4472 not 4298(1867) ; 4298(1867)*
g4473 not 4299(1912) ; 4299(1912)*
g4474 not 7291(1868) ; 7291(1868)*
g4475 not 7292(1881) ; 7292(1881)*
g4476 not 3543(1869) ; 3543(1869)*
g4477 not 3544(1922) ; 3544(1922)*
g4478 not 3091(1870) ; 3091(1870)*
g4479 not 3092(1888) ; 3092(1888)*
g4480 not 4196(1605) ; 4196(1605)*
g4481 not 4197(1921) ; 4197(1921)*
g4482 not 3120(1871) ; 3120(1871)*
g4483 not 3121(1894) ; 3121(1894)*
g4484 not 4178(1872) ; 4178(1872)*
g4485 not 4179(1608) ; 4179(1608)*
g4486 not 3525(1873) ; 3525(1873)*
g4487 not 3526(1610) ; 3526(1610)*
g4488 not 4315(1877) ; 4315(1877)*
g4489 not 4316(1899) ; 4316(1899)*
g4490 not 4219(1942) ; 4219(1942)*
g4491 not 4220(1619) ; 4220(1619)*
g4492 not 3566(1940) ; 3566(1940)*
g4493 not 3567(1878) ; 3567(1878)*
g4494 not 4289(1880) ; 4289(1880)*
g4495 not 4290(1911) ; 4290(1911)*
g4496 not 3534(1882) ; 3534(1882)*
g4497 not 3535(1885) ; 3535(1885)*
g4498 not 3108(1883) ; 3108(1883)*
g4499 not 3109(1892) ; 3109(1892)*
g4500 not 4187(1884) ; 4187(1884)*
g4501 not 4188(1887) ; 4188(1887)*
g4502 not 3100(1886) ; 3100(1886)*
g4503 not 3101(1907) ; 3101(1907)*
g4504 not 4593(1889) ; 4593(1889)*
g4505 not 4594(1890) ; 4594(1890)*
g4506 not 3080(1920) ; 3080(1920)*
g4507 not 3081(1641) ; 3081(1641)*
g4508 not 3117(1930) ; 3117(1930)*
g4509 not 3118(1644) ; 3118(1644)*
g4510 not 7583(1891) ; 7583(1891)*
g4511 not 7584(1906) ; 7584(1906)*
g4512 not 4584(1893) ; 4584(1893)*
g4513 not 4585(1908) ; 4585(1908)*
g4514 not 4575(1909) ; 4575(1909)*
g4515 not 4576(1650) ; 4576(1650)*
g4516 not 4561(1897) ; 4561(1897)*
g4517 not 4562(1895) ; 4562(1895)*
g4518 not 4334(1939) ; 4334(1939)*
g4519 not 4335(1653) ; 4335(1653)*
g4520 not 4325(1941) ; 4325(1941)*
g4521 not 4326(1655) ; 4326(1655)*
g4522 not 4570(1896) ; 4570(1896)*
g4523 not 4571(1898) ; 4571(1898)*
g4524 not 4342(1936) ; 4342(1936)*
g4525 not 4343(1658) ; 4343(1658)*
g4526 not 6763(1918) ; 6763(1918)*
g4527 not 6764(1901) ; 6764(1901)*
g4528 not 3050(1903) ; 3050(1903)*
g4529 not 3051(1669) ; 3051(1669)*
g4530 not 7593(1905) ; 7593(1905)*
g4531 not 7594(1904) ; 7594(1904)*
g4532 not 3060(1919) ; 3060(1919)*
g4533 not 3061(1672) ; 3061(1672)*
g4534 not 3069(1934) ; 3069(1934)*
g4535 not 3070(1675) ; 3070(1675)*
g4536 not 7549(1913) ; 7549(1913)*
g4537 not 7550(1910) ; 7550(1910)*
g4538 not 7539(1916) ; 7539(1916)*
g4539 not 7540(1914) ; 7540(1914)*
g4540 not 3548(1924) ; 3548(1924)*
g4541 not 3549(1696) ; 3549(1696)*
g4542 not 4970(718) ; 4970(718)*
g4543 not 4977(1835) ; 4977(1835)*
g4544 not 4929(564) ; 4929(564)*
g4545 not 4936(1834) ; 4936(1834)*
g4546 not 6753(1932) ; 6753(1932)*
g4547 not 6754(1933) ; 6754(1933)*
g4548 not 3557(1935) ; 3557(1935)*
g4549 not 3558(1938) ; 3558(1938)*
g4550 not 4353(1720) ; 4353(1720)*
g4551 not 4354(1943) ; 4354(1943)*
g4552 not 5929(1048) ; 5929(1048)*
g4553 not 5936(1949) ; 5936(1949)*
g4554 not 6049(1049) ; 6049(1049)*
g4555 not 6056(1948) ; 6056(1948)*
g4556 not 7595(1801) ; 7595(1801)*
g4557 not 7602(2021) ; 7602(2021)*
g4558 not 1816(875) ; 1816(875)*
g4559 not 1945(2019) ; 1945(2019)*
g4560 not 1946(2033) ; 1946(2033)*
g4561 not 1567(876) ; 1567(876)*
g4562 not 1712(2014) ; 1712(2014)*
g4563 not 1713(2030) ; 1713(2030)*
g4564 not 1834(878) ; 1834(878)*
g4565 not 1949(2036) ; 1949(2036)*
g4566 not 7598(1809) ; 7598(1809)*
g4567 not 7601(1997) ; 7601(1997)*
g4568 not 5860(2025) ; 5860(2025)*
g4569 not 5863(1520) ; 5863(1520)*
g4570 not 5852(2026) ; 5852(2026)*
g4571 not 5855(1161) ; 5855(1161)*
g4572 not 1624(894) ; 1624(894)*
g4573 not 1737(2056) ; 1737(2056)*
g4574 not 1738(2067) ; 1738(2067)*
g4575 not 1739(2082) ; 1739(2082)*
g4576 not 1647(899) ; 1647(899)*
g4577 not 1743(2070) ; 1743(2070)*
g4578 not 1744(2085) ; 1744(2085)*
g4579 not 821(929) ; 821(929)*
g4580 not 941(2161) ; 941(2161)*
g4581 not 942(2110) ; 942(2110)*
g4582 not 943(2127) ; 943(2127)*
g4583 not 845(980) ; 845(980)*
g4584 not 947(2113) ; 947(2113)*
g4585 not 948(2130) ; 948(2130)*
g4586 not 7337(1902) ; 7337(1902)*
g4587 not 7344(2203) ; 7344(2203)*
g4588 not 4978(1926) ; 4978(1926)*
g4589 not 4979(2200) ; 4979(2200)*
g4590 not 4937(1929) ; 4937(1929)*
g4591 not 4938(2202) ; 4938(2202)*
g4592 not 7340(1931) ; 7340(1931)*
g4593 not 7343(2191) ; 7343(2191)*
g4594 not 2470(1945) ; 2470(1945)*
g4595 not 2471(2209) ; 2471(2209)*
g4596 not 2740(1947) ; 2740(1947)*
g4597 not 2741(2210) ; 2741(2210)*
g4598 not 7353(1954) ; 7353(1954)*
g4599 not 7360(2216) ; 7360(2216)*
g4600 not 7356(1955) ; 7356(1955)*
g4601 not 7359(2215) ; 7359(2215)*
g4602 not 5362(1956) ; 5362(1956)*
g4603 not 5365(2218) ; 5365(2218)*
g4604 not 5359(1957) ; 5359(1957)*
g4605 not 5366(2217) ; 5366(2217)*
g4606 not 3308(1109) ; 3308(1109)*
g4607 not 3441(2240) ; 3441(2240)*
g4608 not 3442(2251) ; 3442(2251)*
g4609 not 3868(1110) ; 3868(1110)*
g4610 not 4014(2241) ; 4014(2241)*
g4611 not 4015(2257) ; 4015(2257)*
g4612 not 3327(1111) ; 3327(1111)*
g4613 not 3445(2254) ; 3445(2254)*
g4614 not 6682(2244) ; 6682(2244)*
g4615 not 6685(1768) ; 6685(1768)*
g4616 not 6674(2245) ; 6674(2245)*
g4617 not 6677(1474) ; 6677(1474)*
g4618 not 3926(1120) ; 3926(1120)*
g4619 not 4039(2275) ; 4039(2275)*
g4620 not 4040(2285) ; 4040(2285)*
g4621 not 4041(2300) ; 4041(2300)*
g4622 not 3949(1122) ; 3949(1122)*
g4623 not 4045(2288) ; 4045(2288)*
g4624 not 4046(2303) ; 4046(2303)*
g4625 not 2366(1130) ; 2366(1130)*
g4626 not 2503(2323) ; 2503(2323)*
g4627 not 2504(2334) ; 2504(2334)*
g4628 not 2612(1131) ; 2612(1131)*
g4629 not 2765(2324) ; 2765(2324)*
g4630 not 2766(2340) ; 2766(2340)*
g4631 not 2384(1132) ; 2384(1132)*
g4632 not 2507(2337) ; 2507(2337)*
g4633 not 5980(2330) ; 5980(2330)*
g4634 not 5983(1789) ; 5983(1789)*
g4635 not 5972(2331) ; 5972(2331)*
g4636 not 5975(1498) ; 5975(1498)*
g4637 not 2670(1141) ; 2670(1141)*
g4638 not 2792(2355) ; 2792(2355)*
g4639 not 2793(2364) ; 2793(2364)*
g4640 not 2794(2528) ; 2794(2528)*
g4641 not 2693(1143) ; 2693(1143)*
g4642 not 2798(2367) ; 2798(2367)*
g4643 not 2799(2531) ; 2799(2531)*
g4644 not 7436(2394) ; 7436(2394)*
g4645 not 7437(2373) ; 7437(2373)*
g4646 not 5817(2384) ; 5817(2384)*
g4647 not 5824(2380) ; 5824(2380)*
g4648 not 5825(2383) ; 5825(2383)*
g4649 not 5832(2381) ; 5832(2381)*
g4650 not 5841(2392) ; 5841(2392)*
g4651 not 5848(2385) ; 5848(2385)*
g4652 not 5833(2393) ; 5833(2393)*
g4653 not 5840(2386) ; 5840(2386)*
g4654 not 5857(1159) ; 5857(1159)*
g4655 not 5864(2397) ; 5864(2397)*
g4656 not 5849(884) ; 5849(884)*
g4657 not 5856(2398) ; 5856(2398)*
g4658 not 5672(2418) ; 5672(2418)*
g4659 not 5675(1541) ; 5675(1541)*
g4660 not 5584(2419) ; 5584(2419)*
g4661 not 5587(1183) ; 5587(1183)*
g4662 not 4980(2511) ; 4980(2511)*
g4663 not 4987(1549) ; 4987(1549)*
g4664 not 4939(2512) ; 4939(2512)*
g4665 not 4946(1837) ; 4946(1837)*
g4666 not 5102(2481) ; 5102(2481)*
g4667 not 5105(1569) ; 5105(1569)*
g4668 not 5014(2482) ; 5014(2482)*
g4669 not 5017(1219) ; 5017(1219)*
g4670 not 7348(2148) ; 7348(2148)*
g4671 not 7351(2471) ; 7351(2471)*
g4672 not 6822(2150) ; 6822(2150)*
g4673 not 6825(2469) ; 6825(2469)*
g4674 not 6819(2152) ; 6819(2152)*
g4675 not 6826(2467) ; 6826(2467)*
g4676 not 7345(2154) ; 7345(2154)*
g4677 not 7352(2464) ; 7352(2464)*
g4678 not 4369(2486) ; 4369(2486)*
g4679 not 89(48) ; 89(48)*
g4680 not 7614(2181) ; 7614(2181)*
g4681 not 7617(2506) ; 7617(2506)*
g4682 not 6809(2190) ; 6809(2190)*
g4683 not 6816(2515) ; 6816(2515)*
g4684 not 6350(2514) ; 6350(2514)*
g4685 not 6351(2505) ; 6351(2505)*
g4686 not 7611(2193) ; 7611(2193)*
g4687 not 7618(2498) ; 7618(2498)*
g4688 not 7603(2196) ; 7603(2196)*
g4689 not 7610(2508) ; 7610(2508)*
g4690 not 7606(2197) ; 7606(2197)*
g4691 not 7609(2507) ; 7609(2507)*
g4692 not 6812(2204) ; 6812(2204)*
g4693 not 6815(2504) ; 6815(2504)*
g4694 not 6340(2539) ; 6340(2539)*
g4695 not 6341(2538) ; 6341(2538)*
g4696 not 5367(2540) ; 5367(2540)*
g4697 not 5368(2541) ; 5368(2541)*
g4698 not 4836(2745) ; 4836(2745)*
g4699 not 4839(316) ; 4839(316)*
g4700 not 2771(2634) ; 2771(2634)*
g4701 not 4526(205) ; 4526(205)*
g4702 not 6639(2560) ; 6639(2560)*
g4703 not 6646(2556) ; 6646(2556)*
g4704 not 6647(2559) ; 6647(2559)*
g4705 not 6654(2557) ; 6654(2557)*
g4706 not 6663(2567) ; 6663(2567)*
g4707 not 6670(2563) ; 6670(2563)*
g4708 not 6655(2568) ; 6655(2568)*
g4709 not 6662(2564) ; 6662(2564)*
g4710 not 6679(1469) ; 6679(1469)*
g4711 not 6686(2570) ; 6686(2570)*
g4712 not 6671(1116) ; 6671(1116)*
g4713 not 6678(2571) ; 6678(2571)*
g4714 not 7132(2589) ; 7132(2589)*
g4715 not 7135(1780) ; 7135(1780)*
g4716 not 7044(2590) ; 7044(2590)*
g4717 not 7047(1485) ; 7047(1485)*
g4718 not 5937(2610) ; 5937(2610)*
g4719 not 5944(2606) ; 5944(2606)*
g4720 not 5945(2609) ; 5945(2609)*
g4721 not 5952(2607) ; 5952(2607)*
g4722 not 5961(2617) ; 5961(2617)*
g4723 not 5968(2613) ; 5968(2613)*
g4724 not 5953(2618) ; 5953(2618)*
g4725 not 5960(2614) ; 5960(2614)*
g4726 not 5977(1493) ; 5977(1493)*
g4727 not 5984(2622) ; 5984(2622)*
g4728 not 5969(1137) ; 5969(1137)*
g4729 not 5976(2623) ; 5976(2623)*
g4730 not 5820(2002) ; 5820(2002)*
g4731 not 5823(2657) ; 5823(2657)*
g4732 not 5828(2003) ; 5828(2003)*
g4733 not 5831(2656) ; 5831(2656)*
g4734 not 5844(2007) ; 5844(2007)*
g4735 not 5847(2663) ; 5847(2663)*
g4736 not 5836(2008) ; 5836(2008)*
g4737 not 5839(2664) ; 5839(2664)*
g4738 not 5526(2662) ; 5526(2662)*
g4739 not 5529(1519) ; 5529(1519)*
g4740 not 2003(2399) ; 2003(2399)*
g4741 not 2004(2666) ; 2004(2666)*
g4742 not 1999(2400) ; 1999(2400)*
g4743 not 2000(2667) ; 2000(2667)*
g4744 not 5468(2665) ; 5468(2665)*
g4745 not 5471(1162) ; 5471(1162)*
g4746 not 4625(2678) ; 4625(2678)*
g4747 not 4626(2404) ; 4626(2404)*
g4748 not 4622(2673) ; 4622(2673)*
g4749 not 4623(2420) ; 4623(2420)*
g4750 not 5669(1182) ; 5669(1182)*
g4751 not 5676(2671) ; 5676(2671)*
g4752 not 5581(911) ; 5581(911)*
g4753 not 5588(2672) ; 5588(2672)*
g4754 not 4983(1191) ; 4983(1191)*
g4755 not 4986(2742) ; 4986(2742)*
g4756 not 4942(1551) ; 4942(1551)*
g4757 not 4945(2743) ; 4945(2743)*
g4758 not 3598(2692) ; 3598(2692)*
g4759 not 3599(2436) ; 3599(2436)*
g4760 not 3595(2688) ; 3595(2688)*
g4761 not 3596(2450) ; 3596(2450)*
g4762 not 5099(1218) ; 5099(1218)*
g4763 not 5106(2712) ; 5106(2712)*
g4764 not 5011(941) ; 5011(941)*
g4765 not 5018(2713) ; 5018(2713)*
g4766 not 4283(2694) ; 4283(2694)*
g4767 not 4284(2456) ; 4284(2456)*
g4768 not 4286(2693) ; 4286(2693)*
g4769 not 4287(2457) ; 4287(2457)*
g4770 not 1320(2696) ; 1320(2696)*
g4771 not 1321(2460) ; 1321(2460)*
g4772 not 1323(2695) ; 1323(2695)*
g4773 not 1324(2461) ; 1324(2461)*
g4774 not 6360(2697) ; 6360(2697)*
g4775 not 6361(2702) ; 6361(2702)*
g4776 not 6827(2700) ; 6827(2700)*
g4777 not 6828(2701) ; 6828(2701)*
g4778 not 7446(2726) ; 7446(2726)*
g4779 not 7447(2735) ; 7447(2735)*
g4780 not 6817(2744) ; 6817(2744)*
g4781 not 6818(2732) ; 6818(2732)*
g4782 not 7456(2737) ; 7456(2737)*
g4783 not 7457(2736) ; 7457(2736)*
g4784 not 6264(2640) ; 6264(2640)*
g4785 not 6267(2208) ; 6267(2208)*
g4786 not 1314(2749) ; 1314(2749)*
g4787 not 1315(2534) ; 1315(2534)*
g4788 not 1317(2748) ; 1317(2748)*
g4789 not 1318(2535) ; 1318(2535)*
g4790 not 1311(2753) ; 1311(2753)*
g4791 not 1312(2542) ; 1312(2542)*
g4792 not 1308(2752) ; 1308(2752)*
g4793 not 1309(2545) ; 1309(2545)*
g4794 not 4833(207) ; 4833(207)*
g4795 not 4840(2879) ; 4840(2879)*
g4796 not 6642(2227) ; 6642(2227)*
g4797 not 6645(2762) ; 6645(2762)*
g4798 not 6650(2228) ; 6650(2228)*
g4799 not 6653(2761) ; 6653(2761)*
g4800 not 6666(2232) ; 6666(2232)*
g4801 not 6669(2767) ; 6669(2767)*
g4802 not 6658(2233) ; 6658(2233)*
g4803 not 6661(2768) ; 6661(2768)*
g4804 not 3487(2574) ; 3487(2574)*
g4805 not 3488(2771) ; 3488(2771)*
g4806 not 6986(2769) ; 6986(2769)*
g4807 not 6989(1769) ; 6989(1769)*
g4808 not 6928(2770) ; 6928(2770)*
g4809 not 6931(1471) ; 6931(1471)*
g4810 not 3483(2577) ; 3483(2577)*
g4811 not 3484(2772) ; 3484(2772)*
g4812 not 7129(1483) ; 7129(1483)*
g4813 not 7136(2776) ; 7136(2776)*
g4814 not 7041(1127) ; 7041(1127)*
g4815 not 7048(2777) ; 7048(2777)*
g4816 not 2761(2783) ; 2761(2783)*
g4817 not 2753(2603) ; 2753(2603)*
g4818 not 5940(2310) ; 5940(2310)*
g4819 not 5943(2791) ; 5943(2791)*
g4820 not 5948(2311) ; 5948(2311)*
g4821 not 5951(2790) ; 5951(2790)*
g4822 not 2499(2782) ; 2499(2782)*
g4823 not 2491(2608) ; 2491(2608)*
g4824 not 5964(2315) ; 5964(2315)*
g4825 not 5967(2796) ; 5967(2796)*
g4826 not 5956(2316) ; 5956(2316)*
g4827 not 5959(2797) ; 5959(2797)*
g4828 not 2559(2624) ; 2559(2624)*
g4829 not 2560(2800) ; 2560(2800)*
g4830 not 6118(2798) ; 6118(2798)*
g4831 not 6121(1790) ; 6121(1790)*
g4832 not 6060(2799) ; 6060(2799)*
g4833 not 6063(1495) ; 6063(1495)*
g4834 not 2555(2627) ; 2555(2627)*
g4835 not 2556(2801) ; 2556(2801)*
g4836 not 4841(2804) ; 4841(2804)*
g4837 not 4848(2631) ; 4848(2631)*
g4838 not 4849(2807) ; 4849(2807)*
g4839 not 4856(2639) ; 4856(2639)*
g4840 not 4857(2810) ; 4857(2810)*
g4841 not 4864(2641) ; 4864(2641)*
g4842 not 4865(2877) ; 4865(2877)*
g4843 not 4872(2649) ; 4872(2649)*
g4844 not 1985(2817) ; 1985(2817)*
g4845 not 1986(2653) ; 1986(2653)*
g4846 not 1988(2818) ; 1988(2818)*
g4847 not 1989(2654) ; 1989(2654)*
g4848 not 1995(2819) ; 1995(2819)*
g4849 not 1996(2658) ; 1996(2658)*
g4850 not 1992(2820) ; 1992(2820)*
g4851 not 1993(2659) ; 1993(2659)*
g4852 not 5523(1158) ; 5523(1158)*
g4853 not 5530(2821) ; 5530(2821)*
g4854 not 5465(885) ; 5465(885)*
g4855 not 5472(2822) ; 5472(2822)*
g4856 not 4627(2827) ; 4627(2827)*
g4857 not 4624(2829) ; 4624(2829)*
g4858 not 5677(2676) ; 5677(2676)*
g4859 not 5678(2832) ; 5678(2832)*
g4860 not 5589(2677) ; 5589(2677)*
g4861 not 5590(2833) ; 5590(2833)*
g4862 not 4988(2834) ; 4988(2834)*
g4863 not 4989(2679) ; 4989(2679)*
g4864 not 4947(2836) ; 4947(2836)*
g4865 not 4948(2680) ; 4948(2680)*
g4866 not 3600(2838) ; 3600(2838)*
g4867 not 3597(2841) ; 3597(2841)*
g4868 not 5107(2690) ; 5107(2690)*
g4869 not 5108(2843) ; 5108(2843)*
g4870 not 5019(2691) ; 5019(2691)*
g4871 not 5020(2844) ; 5020(2844)*
g4872 not 4288(2846) ; 4288(2846)*
g4873 not 4285(2845) ; 4285(2845)*
g4874 not 1325(2848) ; 1325(2848)*
g4875 not 1322(2847) ; 1322(2847)*
g4876 not 4368(2855) ; 4368(2855)*
g4877 not 4360(2699) ; 4360(2699)*
g4878 not 3604(2853) ; 3604(2853)*
g4879 not 3605(2703) ; 3605(2703)*
g4880 not 4274(2852) ; 4274(2852)*
g4881 not 4275(2707) ; 4275(2707)*
g4882 not 4271(2857) ; 4271(2857)*
g4883 not 4272(2710) ; 4272(2710)*
g4884 not 3601(2856) ; 3601(2856)*
g4885 not 3602(2711) ; 3602(2711)*
g4886 not 3610(2873) ; 3610(2873)*
g4887 not 3611(2718) ; 3611(2718)*
g4888 not 4637(2864) ; 4637(2864)*
g4889 not 4638(2723) ; 4638(2723)*
g4890 not 3135(2868) ; 3135(2868)*
g4891 not 3127(2725) ; 3127(2725)*
g4892 not 4634(2863) ; 4634(2863)*
g4893 not 4635(2727) ; 4635(2727)*
g4894 not 4628(2865) ; 4628(2865)*
g4895 not 4629(2730) ; 4629(2730)*
g4896 not 4631(2866) ; 4631(2866)*
g4897 not 4632(2731) ; 4632(2731)*
g4898 not 4277(2876) ; 4277(2876)*
g4899 not 4278(2739) ; 4278(2739)*
g4900 not 4280(2872) ; 4280(2872)*
g4901 not 4281(2740) ; 4281(2740)*
g4902 not 3607(2875) ; 3607(2875)*
g4903 not 3608(2741) ; 3608(2741)*
g4904 not 6261(1944) ; 6261(1944)*
g4905 not 6268(2808) ; 6268(2808)*
g4906 not 6176(2809) ; 6176(2809)*
g4907 not 6179(1946) ; 6179(1946)*
g4908 not 1319(2883) ; 1319(2883)*
g4909 not 1316(2882) ; 1316(2882)*
g4910 not 1313(2886) ; 1313(2886)*
g4911 not 1310(2887) ; 1310(2887)*
g4912 not 3469(2900) ; 3469(2900)*
g4913 not 3470(2758) ; 3470(2758)*
g4914 not 3472(2901) ; 3472(2901)*
g4915 not 3473(2759) ; 3473(2759)*
g4916 not 3479(2902) ; 3479(2902)*
g4917 not 3480(2765) ; 3480(2765)*
g4918 not 3476(2903) ; 3476(2903)*
g4919 not 3477(2766) ; 3477(2766)*
g4920 not 6983(1470) ; 6983(1470)*
g4921 not 6990(2904) ; 6990(2904)*
g4922 not 6925(1115) ; 6925(1115)*
g4923 not 6932(2905) ; 6932(2905)*
g4924 not 7137(2780) ; 7137(2780)*
g4925 not 7138(2913) ; 7138(2913)*
g4926 not 7049(2781) ; 7049(2781)*
g4927 not 7050(2914) ; 7050(2914)*
g4928 not 2541(2918) ; 2541(2918)*
g4929 not 2542(2786) ; 2542(2786)*
g4930 not 2544(2919) ; 2544(2919)*
g4931 not 2545(2787) ; 2545(2787)*
g4932 not 2551(2921) ; 2551(2921)*
g4933 not 2552(2794) ; 2552(2794)*
g4934 not 2548(2922) ; 2548(2922)*
g4935 not 2549(2795) ; 2549(2795)*
g4936 not 6115(1494) ; 6115(1494)*
g4937 not 6122(2923) ; 6122(2923)*
g4938 not 6057(1136) ; 6057(1136)*
g4939 not 6064(2924) ; 6064(2924)*
g4940 not 4844(2345) ; 4844(2345)*
g4941 not 4847(2932) ; 4847(2932)*
g4942 not 4852(2352) ; 4852(2352)*
g4943 not 4855(2935) ; 4855(2935)*
g4944 not 4860(2358) ; 4860(2358)*
g4945 not 4863(2938) ; 4863(2938)*
g4946 not 4868(2371) ; 4868(2371)*
g4947 not 4871(2985) ; 4871(2985)*
g4948 not 7433(2949) ; 7433(2949)*
g4949 not 7442(2814) ; 7442(2814)*
g4950 not 5531(2823) ; 5531(2823)*
g4951 not 5532(2946) ; 5532(2946)*
g4952 not 5473(2826) ; 5473(2826)*
g4953 not 5474(2948) ; 5474(2948)*
g4954 not 5679(2951) ; 5679(2951)*
g4955 not 5686(2830) ; 5686(2830)*
g4956 not 5591(2952) ; 5591(2952)*
g4957 not 5598(2831) ; 5598(2831)*
g4958 not 6829(2957) ; 6829(2957)*
g4959 not 6836(1833) ; 6836(1833)*
g4960 not 4990(2953) ; 4990(2953)*
g4961 not 4997(1555) ; 4997(1555)*
g4962 not 4949(2954) ; 4949(2954)*
g4963 not 4956(1556) ; 4956(1556)*
g4964 not 5109(2959) ; 5109(2959)*
g4965 not 5116(2840) ; 5116(2840)*
g4966 not 5021(2960) ; 5021(2960)*
g4967 not 5028(2842) ; 5028(2842)*
g4968 not 3606(2966) ; 3606(2966)*
g4969 not 3603(2969) ; 3603(2969)*
g4970 not 4276(2967) ; 4276(2967)*
g4971 not 4273(2968) ; 4273(2968)*
g4972 not 3612(2970) ; 3612(2970)*
g4973 not 3609(2984) ; 3609(2984)*
g4974 not 4639(2973) ; 4639(2973)*
g4975 not 4636(2976) ; 4636(2976)*
g4976 not 4633(2978) ; 4633(2978)*
g4977 not 4630(2977) ; 4630(2977)*
g4978 not 4282(2983) ; 4282(2983)*
g4979 not 4279(2982) ; 4279(2982)*
g4980 not 6269(2878) ; 6269(2878)*
g4981 not 6270(2986) ; 6270(2986)*
g4982 not 6173(1723) ; 6173(1723)*
g4983 not 6180(2936) ; 6180(2936)*
g4984 not 5377(2988) ; 5377(2988)*
g4985 not 5384(1953) ; 5384(1953)*
g4986 not 6337(2961) ; 6337(2961)*
g4987 not 6346(2884) ; 6346(2884)*
g4988 not 5385(2962) ; 5385(2962)*
g4989 not 5392(2885) ; 5392(2885)*
g4990 not 5369(2989) ; 5369(2989)*
g4991 not 5376(1961) ; 5376(1961)*
g4992 not 6991(2907) ; 6991(2907)*
g4993 not 6992(3002) ; 6992(3002)*
g4994 not 6933(2908) ; 6933(2908)*
g4995 not 6934(3003) ; 6934(3003)*
g4996 not 7139(3006) ; 7139(3006)*
g4997 not 7146(2911) ; 7146(2911)*
g4998 not 7051(3007) ; 7051(3007)*
g4999 not 7058(2912) ; 7058(2912)*
g5000 not 6123(2926) ; 6123(2926)*
g5001 not 6124(3014) ; 6124(3014)*
g5002 not 6065(2927) ; 6065(2927)*
g5003 not 6066(3015) ; 6066(3015)*
g5004 not 6271(3064) ; 6271(3064)*
g5005 not 6278(2940) ; 6278(2940)*
g5006 not 7438(2650) ; 7438(2650)*
g5007 not 7441(3039) ; 7441(3039)*
g5008 not 5533(3037) ; 5533(3037)*
g5009 not 5540(2660) ; 5540(2660)*
g5010 not 5475(3038) ; 5475(3038)*
g5011 not 5482(2661) ; 5482(2661)*
g5012 not 5682(2674) ; 5682(2674)*
g5013 not 5685(3042) ; 5685(3042)*
g5014 not 5594(2675) ; 5594(2675)*
g5015 not 5597(3043) ; 5597(3043)*
g5016 not 6832(1546) ; 6832(1546)*
g5017 not 6835(3049) ; 6835(3049)*
g5018 not 4993(1203) ; 4993(1203)*
g5019 not 4996(3045) ; 4996(3045)*
g5020 not 4952(1204) ; 4952(1204)*
g5021 not 4955(3046) ; 4955(3046)*
g5022 not 5112(2687) ; 5112(2687)*
g5023 not 5115(3052) ; 5115(3052)*
g5024 not 5024(2689) ; 5024(2689)*
g5025 not 5027(3053) ; 5027(3053)*
g5026 not 6357(3063) ; 6357(3063)*
g5027 not 6366(2963) ; 6366(2963)*
g5028 not 6845(3058) ; 6845(3058)*
g5029 not 6852(2965) ; 6852(2965)*
g5030 not 7443(3061) ; 7443(3061)*
g5031 not 7452(2975) ; 7452(2975)*
g5032 not 6837(3056) ; 6837(3056)*
g5033 not 6844(2979) ; 6844(2979)*
g5034 not 6347(3057) ; 6347(3057)*
g5035 not 6356(2869) ; 6356(2869)*
g5036 not 7453(3062) ; 7453(3062)*
g5037 not 7462(2981) ; 7462(2981)*
g5038 not 6181(2987) ; 6181(2987)*
g5039 not 6182(3065) ; 6182(3065)*
g5040 not 5380(1736) ; 5380(1736)*
g5041 not 5383(3066) ; 5383(3066)*
g5042 not 6342(2750) ; 6342(2750)*
g5043 not 6345(3054) ; 6345(3054)*
g5044 not 5388(2751) ; 5388(2751)*
g5045 not 5391(3055) ; 5391(3055)*
g5046 not 5372(1759) ; 5372(1759)*
g5047 not 5375(3070) ; 5375(3070)*
g5048 not 6993(3076) ; 6993(3076)*
g5049 not 7000(2763) ; 7000(2763)*
g5050 not 6935(3077) ; 6935(3077)*
g5051 not 6942(2764) ; 6942(2764)*
g5052 not 7142(2778) ; 7142(2778)*
g5053 not 7145(3080) ; 7145(3080)*
g5054 not 7054(2779) ; 7054(2779)*
g5055 not 7057(3081) ; 7057(3081)*
g5056 not 6125(3087) ; 6125(3087)*
g5057 not 6132(2792) ; 6132(2792)*
g5058 not 6067(3088) ; 6067(3088)*
g5059 not 6074(2793) ; 6074(2793)*
g5060 not 6183(3131) ; 6183(3131)*
g5061 not 6190(2939) ; 6190(2939)*
g5062 not 6274(2812) ; 6274(2812)*
g5063 not 6277(3130) ; 6277(3130)*
g5064 not 4515(3099) ; 4515(3099)*
g5065 not 4516(3024) ; 4516(3024)*
g5066 not 5536(2387) ; 5536(2387)*
g5067 not 5539(3104) ; 5539(3104)*
g5068 not 5478(2388) ; 5478(2388)*
g5069 not 5481(3105) ; 5481(3105)*
g5070 not 5687(3106) ; 5687(3106)*
g5071 not 5688(3040) ; 5688(3040)*
g5072 not 5599(3107) ; 5599(3107)*
g5073 not 5600(3041) ; 5600(3041)*
g5074 not 3613(3108) ; 3613(3108)*
g5075 not 3614(3044) ; 3614(3044)*
g5076 not 4998(3111) ; 4998(3111)*
g5077 not 4999(3047) ; 4999(3047)*
g5078 not 4957(3112) ; 4957(3112)*
g5079 not 4958(3048) ; 4958(3048)*
g5080 not 3228(2097) ; 3228(2097)*
g5081 not 3242(3098) ; 3242(3098)*
g5082 not 920(2100) ; 920(2100)*
g5083 not 1447(3100) ; 1447(3100)*
g5084 not 5117(3113) ; 5117(3113)*
g5085 not 5118(3050) ; 5118(3050)*
g5086 not 5029(3114) ; 5029(3114)*
g5087 not 5030(3051) ; 5030(3051)*
g5088 not 6362(2849) ; 6362(2849)*
g5089 not 6365(3129) ; 6365(3129)*
g5090 not 6848(2851) ; 6848(2851)*
g5091 not 6851(3120) ; 6851(3120)*
g5092 not 7448(2862) ; 7448(2862)*
g5093 not 7451(3123) ; 7451(3123)*
g5094 not 6840(2867) ; 6840(2867)*
g5095 not 6843(3118) ; 6843(3118)*
g5096 not 6352(2734) ; 6352(2734)*
g5097 not 6355(3119) ; 6355(3119)*
g5098 not 7458(2870) ; 7458(2870)*
g5099 not 7461(3125) ; 7461(3125)*
g5100 not 1329(3132) ; 1329(3132)*
g5101 not 1330(3067) ; 1330(3067)*
g5102 not 2859(3133) ; 2859(3133)*
g5103 not 2860(3068) ; 2860(3068)*
g5104 not 1332(3134) ; 1332(3134)*
g5105 not 1333(3069) ; 1333(3069)*
g5106 not 1326(3135) ; 1326(3135)*
g5107 not 1327(3071) ; 1327(3071)*
g5108 not 6996(2561) ; 6996(2561)*
g5109 not 6999(3140) ; 6999(3140)*
g5110 not 6938(2562) ; 6938(2562)*
g5111 not 6941(3141) ; 6941(3141)*
g5112 not 7147(3142) ; 7147(3142)*
g5113 not 7148(3078) ; 7148(3078)*
g5114 not 7059(3143) ; 7059(3143)*
g5115 not 7060(3079) ; 7060(3079)*
g5116 not 6128(2611) ; 6128(2611)*
g5117 not 6131(3149) ; 6131(3149)*
g5118 not 6070(2612) ; 6070(2612)*
g5119 not 6073(3150) ; 6073(3150)*
g5120 not 6186(2811) ; 6186(2811)*
g5121 not 6189(3187) ; 6189(3187)*
g5122 not 6279(3155) ; 6279(3155)*
g5123 not 6280(3096) ; 6280(3096)*
g5124 not 5541(3159) ; 5541(3159)*
g5125 not 5542(3102) ; 5542(3102)*
g5126 not 5483(3160) ; 5483(3160)*
g5127 not 5484(3103) ; 5484(3103)*
g5128 not 5689(3164) ; 5689(3164)*
g5129 not 5696(2669) ; 5696(2669)*
g5130 not 5601(3166) ; 5601(3166)*
g5131 not 5608(2670) ; 5608(2670)*
g5132 not 4713(3136) ; 4713(3136)*
g5133 not 4720(2430) ; 4720(2430)*
g5134 not 4959(3170) ; 4959(3170)*
g5135 not 4966(1198) ; 4966(1198)*
g5136 not 5000(3169) ; 5000(3169)*
g5137 not 5007(1201) ; 5007(1201)*
g5138 not 5119(3175) ; 5119(3175)*
g5139 not 5126(2685) ; 5126(2685)*
g5140 not 5031(3178) ; 5031(3178)*
g5141 not 5038(2686) ; 5038(2686)*
g5142 not 4753(3158) ; 4753(3158)*
g5143 not 4760(2455) ; 4760(2455)*
g5144 not 2865(3180) ; 2865(3180)*
g5145 not 2866(3115) ; 2866(3115)*
g5146 not 3619(3181) ; 3619(3181)*
g5147 not 3620(3117) ; 3620(3117)*
g5148 not 3136(2475) ; 3136(2475)*
g5149 not 3149(3182) ; 3149(3182)*
g5150 not 4518(3183) ; 4518(3183)*
g5151 not 4519(3124) ; 4519(3124)*
g5152 not 3616(3184) ; 3616(3184)*
g5153 not 3617(3126) ; 3617(3126)*
g5154 not 2862(3185) ; 2862(3185)*
g5155 not 2863(3127) ; 2863(3127)*
g5156 not 4521(3186) ; 4521(3186)*
g5157 not 4522(3128) ; 4522(3128)*
g5158 not 7001(3193) ; 7001(3193)*
g5159 not 7002(3138) ; 7002(3138)*
g5160 not 6943(3194) ; 6943(3194)*
g5161 not 6944(3139) ; 6944(3139)*
g5162 not 7149(3198) ; 7149(3198)*
g5163 not 7156(2774) ; 7156(2774)*
g5164 not 7061(3199) ; 7061(3199)*
g5165 not 7068(2775) ; 7068(2775)*
g5166 not 4793(3203) ; 4793(3203)*
g5167 not 4800(2598) ; 4800(2598)*
g5168 not 6133(3204) ; 6133(3204)*
g5169 not 6134(3146) ; 6134(3146)*
g5170 not 6075(3205) ; 6075(3205)*
g5171 not 6076(3147) ; 6076(3147)*
g5172 not 6281(3209) ; 6281(3209)*
g5173 not 6288(2805) ; 6288(2805)*
g5174 not 6191(3208) ; 6191(3208)*
g5175 not 6192(3154) ; 6192(3154)*
g5176 not 5543(3212) ; 5543(3212)*
g5177 not 5550(2401) ; 5550(2401)*
g5178 not 5485(3213) ; 5485(3213)*
g5179 not 5492(2402) ; 5492(2402)*
g5180 not 4721(3217) ; 4721(3217)*
g5181 not 4728(2412) ; 4728(2412)*
g5182 not 5692(2413) ; 5692(2413)*
g5183 not 5695(3219) ; 5695(3219)*
g5184 not 5604(2414) ; 5604(2414)*
g5185 not 5607(3221) ; 5607(3221)*
g5186 not 4729(3218) ; 4729(3218)*
g5187 not 4736(2415) ; 4736(2415)*
g5188 not 4737(3220) ; 4737(3220)*
g5189 not 4744(2423) ; 4744(2423)*
g5190 not 4745(3222) ; 4745(3222)*
g5191 not 4752(2425) ; 4752(2425)*
g5192 not 4716(2094) ; 4716(2094)*
g5193 not 4719(3192) ; 4719(3192)*
g5194 not 4962(919) ; 4962(919)*
g5195 not 4965(3227) ; 4965(3227)*
g5196 not 5003(920) ; 5003(920)*
g5197 not 5006(3226) ; 5006(3226)*
g5198 not 4761(3233) ; 4761(3233)*
g5199 not 4768(2442) ; 4768(2442)*
g5200 not 5122(2443) ; 5122(2443)*
g5201 not 5125(3234) ; 5125(3234)*
g5202 not 5034(2444) ; 5034(2444)*
g5203 not 5037(3236) ; 5037(3236)*
g5204 not 4769(3242) ; 4769(3242)*
g5205 not 4776(2445) ; 4776(2445)*
g5206 not 4785(3237) ; 4785(3237)*
g5207 not 4792(2449) ; 4792(2449)*
g5208 not 4756(2139) ; 4756(2139)*
g5209 not 4759(3211) ; 4759(3211)*
g5210 not 4777(3235) ; 4777(3235)*
g5211 not 4784(2485) ; 4784(2485)*
g5212 not 7003(3247) ; 7003(3247)*
g5213 not 7010(2575) ; 7010(2575)*
g5214 not 6945(3248) ; 6945(3248)*
g5215 not 6952(2576) ; 6952(2576)*
g5216 not 4801(3250) ; 4801(3250)*
g5217 not 4808(2583) ; 4808(2583)*
g5218 not 7152(2584) ; 7152(2584)*
g5219 not 7155(3255) ; 7155(3255)*
g5220 not 7064(2585) ; 7064(2585)*
g5221 not 7067(3256) ; 7067(3256)*
g5222 not 4809(3253) ; 4809(3253)*
g5223 not 4816(2586) ; 4816(2586)*
g5224 not 4817(3254) ; 4817(3254)*
g5225 not 4824(2593) ; 4824(2593)*
g5226 not 4825(3257) ; 4825(3257)*
g5227 not 4832(2597) ; 4832(2597)*
g5228 not 4796(2304) ; 4796(2304)*
g5229 not 4799(3259) ; 4799(3259)*
g5230 not 6135(3260) ; 6135(3260)*
g5231 not 6142(2625) ; 6142(2625)*
g5232 not 6077(3261) ; 6077(3261)*
g5233 not 6084(2626) ; 6084(2626)*
g5234 not 6284(2635) ; 6284(2635)*
g5235 not 6287(3264) ; 6287(3264)*
g5236 not 6193(3263) ; 6193(3263)*
g5237 not 6200(2933) ; 6200(2933)*
g5238 not 5546(2038) ; 5546(2038)*
g5239 not 5549(3268) ; 5549(3268)*
g5240 not 5488(2039) ; 5488(2039)*
g5241 not 5491(3269) ; 5491(3269)*
g5242 not 4724(2048) ; 4724(2048)*
g5243 not 4727(3278) ; 4727(3278)*
g5244 not 5697(3276) ; 5697(3276)*
g5245 not 5698(3215) ; 5698(3215)*
g5246 not 5609(3277) ; 5609(3277)*
g5247 not 5610(3216) ; 5610(3216)*
g5248 not 4732(2051) ; 4732(2051)*
g5249 not 4735(3280) ; 4735(3280)*
g5250 not 4740(2066) ; 4740(2066)*
g5251 not 4743(3282) ; 4743(3282)*
g5252 not 4748(2075) ; 4748(2075)*
g5253 not 4751(3284) ; 4751(3284)*
g5254 not 4967(3288) ; 4967(3288)*
g5255 not 4968(3224) ; 4968(3224)*
g5256 not 5008(3289) ; 5008(3289)*
g5257 not 5009(3225) ; 5009(3225)*
g5258 not 4764(2102) ; 4764(2102)*
g5259 not 4767(3297) ; 4767(3297)*
g5260 not 5127(3295) ; 5127(3295)*
g5261 not 5128(3231) ; 5128(3231)*
g5262 not 5039(3296) ; 5039(3296)*
g5263 not 5040(3232) ; 5040(3232)*
g5264 not 4772(2105) ; 4772(2105)*
g5265 not 4775(3303) ; 4775(3303)*
g5266 not 4788(2118) ; 4788(2118)*
g5267 not 4791(3301) ; 4791(3301)*
g5268 not 4780(2168) ; 4780(2168)*
g5269 not 4783(3299) ; 4783(3299)*
g5270 not 7006(2259) ; 7006(2259)*
g5271 not 7009(3312) ; 7009(3312)*
g5272 not 6948(2260) ; 6948(2260)*
g5273 not 6951(3313) ; 6951(3313)*
g5274 not 4804(2266) ; 4804(2266)*
g5275 not 4807(3321) ; 4807(3321)*
g5276 not 7157(3322) ; 7157(3322)*
g5277 not 7158(3251) ; 7158(3251)*
g5278 not 7069(3323) ; 7069(3323)*
g5279 not 7070(3252) ; 7070(3252)*
g5280 not 4812(2269) ; 4812(2269)*
g5281 not 4815(3325) ; 4815(3325)*
g5282 not 4820(2281) ; 4820(2281)*
g5283 not 4823(3327) ; 4823(3327)*
g5284 not 4828(2293) ; 4828(2293)*
g5285 not 4831(3329) ; 4831(3329)*
g5286 not 6138(2342) ; 6138(2342)*
g5287 not 6141(3331) ; 6141(3331)*
g5288 not 6080(2343) ; 6080(2343)*
g5289 not 6083(3332) ; 6083(3332)*
g5290 not 6289(3335) ; 6289(3335)*
g5291 not 6290(3262) ; 6290(3262)*
g5292 not 6196(2806) ; 6196(2806)*
g5293 not 6199(3337) ; 6199(3337)*
g5294 not 5551(3344) ; 5551(3344)*
g5295 not 5552(3272) ; 5552(3272)*
g5296 not 5493(3345) ; 5493(3345)*
g5297 not 5494(3273) ; 5494(3273)*
g5298 not 5699(3347) ; 5699(3347)*
g5299 not 5706(2428) ; 5706(2428)*
g5300 not 5611(3348) ; 5611(3348)*
g5301 not 5618(2429) ; 5618(2429)*
g5302 not 5129(3359) ; 5129(3359)*
g5303 not 5136(2453) ; 5136(2453)*
g5304 not 5041(3360) ; 5041(3360)*
g5305 not 5048(2454) ; 5048(2454)*
g5306 not 7011(3373) ; 7011(3373)*
g5307 not 7012(3315) ; 7012(3315)*
g5308 not 6953(3374) ; 6953(3374)*
g5309 not 6954(3316) ; 6954(3316)*
g5310 not 7159(3377) ; 7159(3377)*
g5311 not 7166(2599) ; 7166(2599)*
g5312 not 7071(3378) ; 7071(3378)*
g5313 not 7078(2600) ; 7078(2600)*
g5314 not 6143(3383) ; 6143(3383)*
g5315 not 6144(3333) ; 6144(3333)*
g5316 not 6085(3384) ; 6085(3384)*
g5317 not 6086(3334) ; 6086(3334)*
g5318 not 6201(3386) ; 6201(3386)*
g5319 not 6202(3336) ; 6202(3336)*
g5320 not 5495(3392) ; 5495(3392)*
g5321 not 5502(2395) ; 5502(2395)*
g5322 not 5553(3391) ; 5553(3391)*
g5323 not 5560(2396) ; 5560(2396)*
g5324 not 5702(2090) ; 5702(2090)*
g5325 not 5705(3394) ; 5705(3394)*
g5326 not 5614(2091) ; 5614(2091)*
g5327 not 5617(3395) ; 5617(3395)*
g5328 not 5132(2135) ; 5132(2135)*
g5329 not 5135(3409) ; 5135(3409)*
g5330 not 5044(2136) ; 5044(2136)*
g5331 not 5047(3410) ; 5047(3410)*
g5332 not 6291(3385) ; 6291(3385)*
g5333 not 6298(2880) ; 6298(2880)*
g5334 not 6955(3423) ; 6955(3423)*
g5335 not 6962(2572) ; 6962(2572)*
g5336 not 7013(3422) ; 7013(3422)*
g5337 not 7020(2573) ; 7020(2573)*
g5338 not 7162(2305) ; 7162(2305)*
g5339 not 7165(3427) ; 7165(3427)*
g5340 not 7074(2306) ; 7074(2306)*
g5341 not 7077(3428) ; 7077(3428)*
g5342 not 6087(3435) ; 6087(3435)*
g5343 not 6094(2620) ; 6094(2620)*
g5344 not 6145(3434) ; 6145(3434)*
g5345 not 6152(2621) ; 6152(2621)*
g5346 not 5498(2023) ; 5498(2023)*
g5347 not 5501(3441) ; 5501(3441)*
g5348 not 5556(2024) ; 5556(2024)*
g5349 not 5559(3440) ; 5559(3440)*
g5350 not 5707(3442) ; 5707(3442)*
g5351 not 5708(3399) ; 5708(3399)*
g5352 not 5619(3443) ; 5619(3443)*
g5353 not 5620(3400) ; 5620(3400)*
g5354 not 5137(3447) ; 5137(3447)*
g5355 not 5138(3413) ; 5138(3413)*
g5356 not 5049(3448) ; 5049(3448)*
g5357 not 5050(3414) ; 5050(3414)*
g5358 not 6294(2746) ; 6294(2746)*
g5359 not 6297(3436) ; 6297(3436)*
g5360 not 6203(3437) ; 6203(3437)*
g5361 not 6210(2881) ; 6210(2881)*
g5362 not 6958(2248) ; 6958(2248)*
g5363 not 6961(3457) ; 6961(3457)*
g5364 not 7016(2249) ; 7016(2249)*
g5365 not 7019(3456) ; 7019(3456)*
g5366 not 7167(3458) ; 7167(3458)*
g5367 not 7168(3432) ; 7168(3432)*
g5368 not 7079(3459) ; 7079(3459)*
g5369 not 7080(3433) ; 7080(3433)*
g5370 not 6090(2328) ; 6090(2328)*
g5371 not 6093(3463) ; 6093(3463)*
g5372 not 6148(2329) ; 6148(2329)*
g5373 not 6151(3462) ; 6151(3462)*
g5374 not 5503(3465) ; 5503(3465)*
g5375 not 5504(3438) ; 5504(3438)*
g5376 not 5561(3466) ; 5561(3466)*
g5377 not 5562(3439) ; 5562(3439)*
g5378 not 5621(3468) ; 5621(3468)*
g5379 not 5628(2426) ; 5628(2426)*
g5380 not 5709(3467) ; 5709(3467)*
g5381 not 5716(2427) ; 5716(2427)*
g5382 not 5051(3471) ; 5051(3471)*
g5383 not 5058(2451) ; 5058(2451)*
g5384 not 5139(3470) ; 5139(3470)*
g5385 not 5146(2452) ; 5146(2452)*
g5386 not 6299(3472) ; 6299(3472)*
g5387 not 6300(3453) ; 6300(3453)*
g5388 not 6206(2747) ; 6206(2747)*
g5389 not 6209(3464) ; 6209(3464)*
g5390 not 6963(3474) ; 6963(3474)*
g5391 not 6964(3454) ; 6964(3454)*
g5392 not 7021(3475) ; 7021(3475)*
g5393 not 7022(3455) ; 7022(3455)*
g5394 not 7081(3477) ; 7081(3477)*
g5395 not 7088(2595) ; 7088(2595)*
g5396 not 7169(3476) ; 7169(3476)*
g5397 not 7176(2596) ; 7176(2596)*
g5398 not 6095(3478) ; 6095(3478)*
g5399 not 6096(3460) ; 6096(3460)*
g5400 not 6153(3479) ; 6153(3479)*
g5401 not 6154(3461) ; 6154(3461)*
g5402 not 6301(3490) ; 6301(3490)*
g5403 not 6308(2647) ; 6308(2647)*
g5404 not 5563(3481) ; 5563(3481)*
g5405 not 5570(2376) ; 5570(2376)*
g5406 not 5505(3480) ; 5505(3480)*
g5407 not 5512(2377) ; 5512(2377)*
g5408 not 5624(2076) ; 5624(2076)*
g5409 not 5627(3485) ; 5627(3485)*
g5410 not 5712(2077) ; 5712(2077)*
g5411 not 5715(3484) ; 5715(3484)*
g5412 not 5054(2121) ; 5054(2121)*
g5413 not 5057(3489) ; 5057(3489)*
g5414 not 5142(2123) ; 5142(2123)*
g5415 not 5145(3488) ; 5145(3488)*
g5416 not 6211(3491) ; 6211(3491)*
g5417 not 6212(3473) ; 6212(3473)*
g5418 not 7023(3493) ; 7023(3493)*
g5419 not 7030(2554) ; 7030(2554)*
g5420 not 6965(3492) ; 6965(3492)*
g5421 not 6972(2555) ; 6972(2555)*
g5422 not 7084(2290) ; 7084(2290)*
g5423 not 7087(3497) ; 7087(3497)*
g5424 not 7172(2291) ; 7172(2291)*
g5425 not 7175(3496) ; 7175(3496)*
g5426 not 6155(3499) ; 6155(3499)*
g5427 not 6162(2604) ; 6162(2604)*
g5428 not 6097(3498) ; 6097(3498)*
g5429 not 6104(2605) ; 6104(2605)*
g5430 not 6213(3510) ; 6213(3510)*
g5431 not 6220(2646) ; 6220(2646)*
g5432 not 6304(2370) ; 6304(2370)*
g5433 not 6307(3509) ; 6307(3509)*
g5434 not 5566(2000) ; 5566(2000)*
g5435 not 5569(3504) ; 5569(3504)*
g5436 not 5508(2001) ; 5508(2001)*
g5437 not 5511(3503) ; 5511(3503)*
g5438 not 5629(3505) ; 5629(3505)*
g5439 not 5630(3482) ; 5630(3482)*
g5440 not 5717(3506) ; 5717(3506)*
g5441 not 5718(3483) ; 5718(3483)*
g5442 not 5059(3507) ; 5059(3507)*
g5443 not 5060(3486) ; 5060(3486)*
g5444 not 5147(3508) ; 5147(3508)*
g5445 not 5148(3487) ; 5148(3487)*
g5446 not 7026(2225) ; 7026(2225)*
g5447 not 7029(3514) ; 7029(3514)*
g5448 not 6968(2226) ; 6968(2226)*
g5449 not 6971(3513) ; 6971(3513)*
g5450 not 7089(3515) ; 7089(3515)*
g5451 not 7090(3494) ; 7090(3494)*
g5452 not 7177(3516) ; 7177(3516)*
g5453 not 7178(3495) ; 7178(3495)*
g5454 not 6158(2308) ; 6158(2308)*
g5455 not 6161(3520) ; 6161(3520)*
g5456 not 6100(2309) ; 6100(2309)*
g5457 not 6103(3519) ; 6103(3519)*
g5458 not 6216(2369) ; 6216(2369)*
g5459 not 6219(3529) ; 6219(3529)*
g5460 not 6309(3522) ; 6309(3522)*
g5461 not 6310(3500) ; 6310(3500)*
g5462 not 5571(3523) ; 5571(3523)*
g5463 not 5572(3501) ; 5572(3501)*
g5464 not 5513(3524) ; 5513(3524)*
g5465 not 5514(3502) ; 5514(3502)*
g5466 not 5719(3526) ; 5719(3526)*
g5467 not 5726(2408) ; 5726(2408)*
g5468 not 5631(3525) ; 5631(3525)*
g5469 not 5638(2409) ; 5638(2409)*
g5470 not 5149(3528) ; 5149(3528)*
g5471 not 5156(2439) ; 5156(2439)*
g5472 not 5061(3527) ; 5061(3527)*
g5473 not 5068(2440) ; 5068(2440)*
g5474 not 7031(3530) ; 7031(3530)*
g5475 not 7032(3511) ; 7032(3511)*
g5476 not 6973(3531) ; 6973(3531)*
g5477 not 6974(3512) ; 6974(3512)*
g5478 not 7179(3533) ; 7179(3533)*
g5479 not 7186(2580) ; 7186(2580)*
g5480 not 7091(3532) ; 7091(3532)*
g5481 not 7098(2581) ; 7098(2581)*
g5482 not 6163(3534) ; 6163(3534)*
g5483 not 6164(3517) ; 6164(3517)*
g5484 not 6105(3535) ; 6105(3535)*
g5485 not 6106(3518) ; 6106(3518)*
g5486 not 6311(3537) ; 6311(3537)*
g5487 not 6318(2632) ; 6318(2632)*
g5488 not 6221(3536) ; 6221(3536)*
g5489 not 6222(3521) ; 6222(3521)*
g5490 not 5515(3539) ; 5515(3539)*
g5491 not 5522(2389) ; 5522(2389)*
g5492 not 5573(3538) ; 5573(3538)*
g5493 not 5580(2390) ; 5580(2390)*
g5494 not 5722(2044) ; 5722(2044)*
g5495 not 5725(3543) ; 5725(3543)*
g5496 not 5634(2045) ; 5634(2045)*
g5497 not 5637(3542) ; 5637(3542)*
g5498 not 5152(2098) ; 5152(2098)*
g5499 not 5155(3547) ; 5155(3547)*
g5500 not 5064(2099) ; 5064(2099)*
g5501 not 5067(3546) ; 5067(3546)*
g5502 not 6975(3549) ; 6975(3549)*
g5503 not 6982(2565) ; 6982(2565)*
g5504 not 7033(3548) ; 7033(3548)*
g5505 not 7040(2566) ; 7040(2566)*
g5506 not 7182(2262) ; 7182(2262)*
g5507 not 7185(3553) ; 7185(3553)*
g5508 not 7094(2263) ; 7094(2263)*
g5509 not 7097(3552) ; 7097(3552)*
g5510 not 6107(3555) ; 6107(3555)*
g5511 not 6114(2615) ; 6114(2615)*
g5512 not 6165(3554) ; 6165(3554)*
g5513 not 6172(2616) ; 6172(2616)*
g5514 not 6314(2346) ; 6314(2346)*
g5515 not 6317(3558) ; 6317(3558)*
g5516 not 6223(3557) ; 6223(3557)*
g5517 not 6230(2633) ; 6230(2633)*
g5518 not 5518(2011) ; 5518(2011)*
g5519 not 5521(3560) ; 5521(3560)*
g5520 not 5576(2013) ; 5576(2013)*
g5521 not 5579(3559) ; 5579(3559)*
g5522 not 5727(3563) ; 5727(3563)*
g5523 not 5728(3540) ; 5728(3540)*
g5524 not 5639(3564) ; 5639(3564)*
g5525 not 5640(3541) ; 5640(3541)*
g5526 not 5157(3565) ; 5157(3565)*
g5527 not 5158(3544) ; 5158(3544)*
g5528 not 5069(3566) ; 5069(3566)*
g5529 not 5070(3545) ; 5070(3545)*
g5530 not 6978(2235) ; 6978(2235)*
g5531 not 6981(3568) ; 6981(3568)*
g5532 not 7036(2237) ; 7036(2237)*
g5533 not 7039(3567) ; 7039(3567)*
g5534 not 7187(3571) ; 7187(3571)*
g5535 not 7188(3550) ; 7188(3550)*
g5536 not 7099(3572) ; 7099(3572)*
g5537 not 7100(3551) ; 7100(3551)*
g5538 not 6110(2318) ; 6110(2318)*
g5539 not 6113(3574) ; 6113(3574)*
g5540 not 6168(2320) ; 6168(2320)*
g5541 not 6171(3573) ; 6171(3573)*
g5542 not 6319(3577) ; 6319(3577)*
g5543 not 6320(3556) ; 6320(3556)*
g5544 not 6226(2347) ; 6226(2347)*
g5545 not 6229(3579) ; 6229(3579)*
g5546 not 1755(3580) ; 1755(3580)*
g5547 not 1756(3561) ; 1756(3561)*
g5548 not 1760(3581) ; 1760(3581)*
g5549 not 1761(3562) ; 1761(3562)*
g5550 not 5729(3582) ; 5729(3582)*
g5551 not 5736(2421) ; 5736(2421)*
g5552 not 5641(3583) ; 5641(3583)*
g5553 not 5648(2422) ; 5648(2422)*
g5554 not 5159(3584) ; 5159(3584)*
g5555 not 5166(2483) ; 5166(2483)*
g5556 not 5071(3585) ; 5071(3585)*
g5557 not 5078(2484) ; 5078(2484)*
g5558 not 4057(3586) ; 4057(3586)*
g5559 not 4058(3569) ; 4058(3569)*
g5560 not 4062(3587) ; 4062(3587)*
g5561 not 4063(3570) ; 4063(3570)*
g5562 not 7189(3588) ; 7189(3588)*
g5563 not 7196(2591) ; 7196(2591)*
g5564 not 7101(3589) ; 7101(3589)*
g5565 not 7108(2592) ; 7108(2592)*
g5566 not 2817(3590) ; 2817(3590)*
g5567 not 2818(3575) ; 2818(3575)*
g5568 not 2822(3591) ; 2822(3591)*
g5569 not 2823(3576) ; 2823(3576)*
g5570 not 6231(3593) ; 6231(3593)*
g5571 not 6232(3578) ; 6232(3578)*
g5572 not 6321(3592) ; 6321(3592)*
g5573 not 6328(2642) ; 6328(2642)*
g5574 not 5732(2063) ; 5732(2063)*
g5575 not 5735(3596) ; 5735(3596)*
g5576 not 5644(2064) ; 5644(2064)*
g5577 not 5647(3597) ; 5647(3597)*
g5578 not 5162(2166) ; 5162(2166)*
g5579 not 5165(3600) ; 5165(3600)*
g5580 not 5074(2167) ; 5074(2167)*
g5581 not 5077(3601) ; 5077(3601)*
g5582 not 7192(2278) ; 7192(2278)*
g5583 not 7195(3606) ; 7195(3606)*
g5584 not 7104(2279) ; 7104(2279)*
g5585 not 7107(3607) ; 7107(3607)*
g5586 not 6324(2359) ; 6324(2359)*
g5587 not 6327(3612) ; 6327(3612)*
g5588 not 6233(3613) ; 6233(3613)*
g5589 not 6240(2643) ; 6240(2643)*
g5590 not 5659(3619) ; 5659(3619)*
g5591 not 5660(3598) ; 5660(3598)*
g5592 not 5649(3620) ; 5649(3620)*
g5593 not 5650(3599) ; 5650(3599)*
g5594 not 5089(3621) ; 5089(3621)*
g5595 not 5090(3602) ; 5090(3602)*
g5596 not 5079(3622) ; 5079(3622)*
g5597 not 5080(3603) ; 5080(3603)*
g5598 not 7119(3631) ; 7119(3631)*
g5599 not 7120(3608) ; 7120(3608)*
g5600 not 7109(3632) ; 7109(3632)*
g5601 not 7110(3609) ; 7110(3609)*
g5602 not 6251(3634) ; 6251(3634)*
g5603 not 6252(3614) ; 6252(3614)*
g5604 not 6236(2360) ; 6236(2360)*
g5605 not 6239(3633) ; 6239(3633)*
g5606 not 5661(3637) ; 5661(3637)*
g5607 not 5668(2416) ; 5668(2416)*
g5608 not 5651(3638) ; 5651(3638)*
g5609 not 5658(2417) ; 5658(2417)*
g5610 not 5091(3639) ; 5091(3639)*
g5611 not 5098(2446) ; 5098(2446)*
g5612 not 5081(3640) ; 5081(3640)*
g5613 not 5088(2447) ; 5088(2447)*
g5614 not 7121(3643) ; 7121(3643)*
g5615 not 7128(2587) ; 7128(2587)*
g5616 not 7111(3644) ; 7111(3644)*
g5617 not 7118(2588) ; 7118(2588)*
g5618 not 6253(3645) ; 6253(3645)*
g5619 not 6260(2636) ; 6260(2636)*
g5620 not 6241(3646) ; 6241(3646)*
g5621 not 6242(3635) ; 6242(3635)*
g5622 not 5664(2052) ; 5664(2052)*
g5623 not 5667(3650) ; 5667(3650)*
g5624 not 5654(2054) ; 5654(2054)*
g5625 not 5657(3651) ; 5657(3651)*
g5626 not 5094(2106) ; 5094(2106)*
g5627 not 5097(3654) ; 5097(3654)*
g5628 not 5084(2108) ; 5084(2108)*
g5629 not 5087(3655) ; 5087(3655)*
g5630 not 7124(2270) ; 7124(2270)*
g5631 not 7127(3660) ; 7127(3660)*
g5632 not 7114(2272) ; 7114(2272)*
g5633 not 7117(3661) ; 7117(3661)*
g5634 not 6256(2350) ; 6256(2350)*
g5635 not 6259(3663) ; 6259(3663)*
g5636 not 6243(3664) ; 6243(3664)*
g5637 not 6250(2638) ; 6250(2638)*
g5638 not 1778(3665) ; 1778(3665)*
g5639 not 1779(3648) ; 1779(3648)*
g5640 not 1775(3666) ; 1775(3666)*
g5641 not 1776(3649) ; 1776(3649)*
g5642 not 987(3667) ; 987(3667)*
g5643 not 988(3652) ; 988(3652)*
g5644 not 984(3668) ; 984(3668)*
g5645 not 985(3653) ; 985(3653)*
g5646 not 4079(3669) ; 4079(3669)*
g5647 not 4080(3658) ; 4080(3658)*
g5648 not 4076(3670) ; 4076(3670)*
g5649 not 4077(3659) ; 4077(3659)*
g5650 not 2840(3671) ; 2840(3671)*
g5651 not 2841(3662) ; 2841(3662)*
g5652 not 6246(2351) ; 6246(2351)*
g5653 not 6249(3673) ; 6249(3673)*
g5654 not 2837(3682) ; 2837(3682)*
g5655 not 2838(3672) ; 2838(3672)*
g5656 not 5740(3694) ; 5740(3694)*
g5657 not 5743(3647) ; 5743(3647)*
g5658 not 5170(3696) ; 5170(3696)*
g5659 not 5173(3469) ; 5173(3469)*
g5660 not 6332(3697) ; 6332(3697)*
g5661 not 6335(3656) ; 6335(3656)*
g5662 not 7200(3699) ; 7200(3699)*
g5663 not 7203(3657) ; 7203(3657)*
g5664 not 5737(3636) ; 5737(3636)*
g5665 not 5744(3698) ; 5744(3698)*
g5666 not 5167(3446) ; 5167(3446)*
g5667 not 5174(3700) ; 5174(3700)*
g5668 not 6329(3641) ; 6329(3641)*
g5669 not 6336(3704) ; 6336(3704)*
g5670 not 7197(3642) ; 7197(3642)*
g5671 not 7204(3706) ; 7204(3706)*
g5672 not 1791(3701) ; 1791(3701)*
g5673 not 1792(3707) ; 1792(3707)*
g5674 not 1003(3702) ; 1003(3702)*
g5675 not 1004(3708) ; 1004(3708)*
g5676 not 2855(3703) ; 2855(3703)*
g5677 not 2856(3709) ; 2856(3709)*
g5678 not 4092(3705) ; 4092(3705)*
g5679 not 4093(3710) ; 4093(3710)*
