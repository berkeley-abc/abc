name C880.iscas
i 1GAT(0)
i 8GAT(1)
i 13GAT(2)
i 17GAT(3)
i 26GAT(4)
i 29GAT(5)
i 36GAT(6)
i 42GAT(7)
i 51GAT(8)
i 55GAT(9)
i 59GAT(10)
i 68GAT(11)
i 72GAT(12)
i 73GAT(13)
i 74GAT(14)
i 75GAT(15)
i 80GAT(16)
i 85GAT(17)
i 86GAT(18)
i 87GAT(19)
i 88GAT(20)
i 89GAT(21)
i 90GAT(22)
i 91GAT(23)
i 96GAT(24)
i 101GAT(25)
i 106GAT(26)
i 111GAT(27)
i 116GAT(28)
i 121GAT(29)
i 126GAT(30)
i 130GAT(31)
i 135GAT(32)
i 138GAT(33)
i 143GAT(34)
i 146GAT(35)
i 149GAT(36)
i 152GAT(37)
i 153GAT(38)
i 156GAT(39)
i 159GAT(40)
i 165GAT(41)
i 171GAT(42)
i 177GAT(43)
i 183GAT(44)
i 189GAT(45)
i 195GAT(46)
i 201GAT(47)
i 207GAT(48)
i 210GAT(49)
i 219GAT(50)
i 228GAT(51)
i 237GAT(52)
i 246GAT(53)
i 255GAT(54)
i 259GAT(55)
i 260GAT(56)
i 261GAT(57)
i 267GAT(58)
i 268GAT(59)

o 388GAT(133)
o 389GAT(132)
o 390GAT(131)
o 391GAT(124)
o 418GAT(168)
o 419GAT(164)
o 420GAT(158)
o 421GAT(162)
o 422GAT(161)
o 423GAT(155)
o 446GAT(183)
o 447GAT(182)
o 448GAT(179)
o 449GAT(176)
o 450GAT(173)
o 767GAT(349)
o 768GAT(334)
o 850GAT(404)
o 863GAT(424)
o 864GAT(423)
o 865GAT(422)
o 866GAT(426)
o 874GAT(433)
o 878GAT(442)
o 879GAT(441)
o 880GAT(440)

g1 and 268GAT(59) ; 310GAT(60)
g2 and 267GAT(58) 255GAT(54) ; 341GAT(61)
g3 and 260GAT(56) 255GAT(54) ; 339GAT(62)
g4 and 259GAT(55) 255GAT(54) ; 337GAT(63)
g5 and 201GAT(47)* 195GAT(46)* ; 331GAT(64)
g6 and 201GAT(47) 195GAT(46) ; 330GAT(65)
g7 and 189GAT(45)* 183GAT(44)* ; 329GAT(66)
g8 and 189GAT(45) 183GAT(44) ; 328GAT(67)
g9 and 177GAT(43)* 171GAT(42)* ; 327GAT(68)
g10 and 177GAT(43) 171GAT(42) ; 326GAT(69)
g11 and 165GAT(41)* 159GAT(40)* ; 325GAT(70)
g12 and 165GAT(41) 159GAT(40) ; 324GAT(71)
g13 and 138GAT(33) 152GAT(37) ; 318GAT(72)
g14 and 121GAT(29) 210GAT(49) ; 340GAT(73)
g15 and 126GAT(30)* 121GAT(29)* ; 308GAT(74)
g16 and 126GAT(30) 121GAT(29) ; 307GAT(75)
g17 and 116GAT(28) 210GAT(49) ; 338GAT(76)
g18 and 111GAT(27) 210GAT(49) ; 336GAT(77)
g19 and 116GAT(28)* 111GAT(27)* ; 306GAT(78)
g20 and 116GAT(28) 111GAT(27) ; 305GAT(79)
g21 and 106GAT(26) 210GAT(49) ; 335GAT(80)
g22 and 101GAT(25) 210GAT(49) ; 334GAT(81)
g23 and 106GAT(26)* 101GAT(25)* ; 304GAT(82)
g24 and 106GAT(26) 101GAT(25) ; 303GAT(83)
g25 and 96GAT(24) 210GAT(49) ; 333GAT(84)
g26 and 91GAT(23) 210GAT(49) ; 332GAT(85)
g27 and 96GAT(24)* 91GAT(23)* ; 302GAT(86)
g28 and 96GAT(24) 91GAT(23) ; 301GAT(87)
g29 and 88GAT(20)* 87GAT(19)* ; 298GAT(88)
g30 and 86GAT(18) 85GAT(17) ; 297GAT(89)
g31 and 156GAT(39) 59GAT(10) ; 319GAT(90)
g32 and 80GAT(16) 75GAT(15) 59GAT(10) ; 293GAT(91)
g33 and 74GAT(14) 68GAT(11) 59GAT(10) ; 286GAT(92)
g34 and 138GAT(33) 51GAT(8) ; 316GAT(93)
g35 and 42GAT(7) 75GAT(15) 59GAT(10) ; 294GAT(94)
g36 and 72GAT(12) 68GAT(11) 42GAT(7) 59GAT(10) ; 284GAT(95)
g37 and 42GAT(7) 36GAT(6) 59GAT(10) ; 296GAT(96)
g38 and 80GAT(16) 36GAT(6) 59GAT(10) ; 295GAT(97)
g39 and 42GAT(7) 36GAT(6) 29GAT(5) ; 292GAT(98)
g40 and 80GAT(16) 36GAT(6) 29GAT(5) ; 291GAT(99)
g41 and 42GAT(7) 75GAT(15) 29GAT(5) ; 290GAT(100)
g42 and 80GAT(16) 75GAT(15) 29GAT(5) ; 287GAT(101)
g43 and 68GAT(11) 29GAT(5) ; 285GAT(102)
g44 and 42GAT(7) 36GAT(6) 29GAT(5) ; 273GAT(103)
g45 and 42GAT(7) 17GAT(3) ; 323GAT(104)
g46 and 42GAT(7)* 17GAT(3)* ; 322GAT(105)
g47 and 138GAT(33) 17GAT(3) ; 317GAT(106)
g48 and 138GAT(33) 8GAT(1) ; 309GAT(107)
g49 and 55GAT(9) 13GAT(2) 8GAT(1) 1GAT(0) ; 280GAT(108)
g50 and 17GAT(3) 51GAT(8) 8GAT(1) 1GAT(0) ; 279GAT(109)
g51 and 51GAT(8) 26GAT(4) 1GAT(0) ; 276GAT(110)
g52 and 17GAT(3) 13GAT(2) 26GAT(4) 1GAT(0) ; 270GAT(111)
g53 and 17GAT(3) 13GAT(2) 8GAT(1) 1GAT(0) ; 269GAT(112)
g54 and 310GAT(60) ; 369GAT(113)
g55 and 331GAT(64) 330GAT(65) ; 385GAT(114)
g56 and 329GAT(66) 328GAT(67) ; 382GAT(115)
g57 and 327GAT(68) 326GAT(69) ; 379GAT(116)
g58 and 325GAT(70) 324GAT(71) ; 376GAT(117)
g59 and 308GAT(74) 307GAT(75) ; 366GAT(118)
g60 and 306GAT(78) 305GAT(79) ; 363GAT(119)
g61 and 304GAT(82) 303GAT(83) ; 360GAT(120)
g62 and 302GAT(86) 301GAT(87) ; 357GAT(121)
g63 and 298GAT(88) 90GAT(22) ; 356GAT(122)
g64 and 298GAT(88) 89GAT(21) ; 355GAT(123)
g65 and 297GAT(89) ; 391GAT(124)
g66 and 293GAT(91) ; 351GAT(125)
g67 and 286GAT(92)* 280GAT(108)* ; 350GAT(126)
g68 and 294GAT(94) ; 352GAT(127)
g69 and 284GAT(95)* 280GAT(108)* ; 348GAT(128)
g70 and 296GAT(96) ; 354GAT(129)
g71 and 295GAT(97) ; 353GAT(130)
g72 and 292GAT(98) ; 390GAT(131)
g73 and 291GAT(99) ; 389GAT(132)
g74 and 290GAT(100) ; 388GAT(133)
g75 and 285GAT(102)* 280GAT(108)* ; 349GAT(134)
g76 and 273GAT(103) ; 343GAT(135)
g77 and 273GAT(103)* 270GAT(111)* ; 344GAT(136)
g78 and 323GAT(104)* 322GAT(105)* ; 375GAT(137)
g79 and 279GAT(109) ; 347GAT(138)
g80 and 276GAT(110) ; 345GAT(139)
g81 and 276GAT(110) ; 346GAT(140)
g82 and 269GAT(112) ; 342GAT(141)
g83 and 369GAT(113) 210GAT(49) ; 417GAT(142)
g84 and 385GAT(114) ; 415GAT(143)
g85 and 385GAT(114) 382GAT(115) ; 416GAT(144)
g86 and 382GAT(115) ; 414GAT(145)
g87 and 379GAT(116) ; 412GAT(146)
g88 and 379GAT(116) 376GAT(117) ; 413GAT(147)
g89 and 376GAT(117) ; 411GAT(148)
g90 and 366GAT(118) ; 408GAT(149)
g91 and 366GAT(118) 363GAT(119) ; 409GAT(150)
g92 and 363GAT(119) ; 407GAT(151)
g93 and 360GAT(120) ; 405GAT(152)
g94 and 360GAT(120) 357GAT(121) ; 406GAT(153)
g95 and 357GAT(121) ; 404GAT(154)
g96 and 356GAT(122) ; 423GAT(155)
g97 and 355GAT(123) ; 403GAT(156)
g98 and 73GAT(13) 348GAT(128) ; 400GAT(157)
g99 and 351GAT(125) ; 420GAT(158)
g100 and 350GAT(126) ; 402GAT(159)
g101 and 352GAT(127) 347GAT(138) ; 410GAT(160)
g102 and 354GAT(129) ; 422GAT(161)
g103 and 353GAT(130) ; 421GAT(162)
g104 and 349GAT(134) ; 401GAT(163)
g105 and 344GAT(136) ; 419GAT(164)
g106 and 345GAT(139) ; 393GAT(165)
g107 and 346GAT(140) ; 399GAT(166)
g108 and 343GAT(135)* 270GAT(111)* ; 392GAT(167)
g109 and 342GAT(141) ; 418GAT(168)
g110 and 415GAT(143) 414GAT(145) ; 445GAT(169)
g111 and 412GAT(146) 411GAT(148) ; 444GAT(170)
g112 and 408GAT(149) 407GAT(151) ; 426GAT(171)
g113 and 405GAT(152) 404GAT(154) ; 425GAT(172)
g114 and 403GAT(156) ; 450GAT(173)
g115 and 400GAT(157) ; 424GAT(174)
g116 and 393GAT(165) 156GAT(39) 59GAT(10) 375GAT(137) ; 442GAT(175)
g117 and 402GAT(159) ; 449GAT(176)
g118 and 55GAT(9) 287GAT(101) 393GAT(165) ; 437GAT(177)
g119 and 55GAT(9) 393GAT(165) 319GAT(90) ; 427GAT(178)
g120 and 401GAT(163) ; 448GAT(179)
g121 and 17GAT(3) 319GAT(90) 393GAT(165) ; 443GAT(180)
g122 and 287GAT(101) 17GAT(3) 393GAT(165) ; 432GAT(181)
g123 and 399GAT(166) ; 447GAT(182)
g124 and 392GAT(167) ; 446GAT(183)
g125 and 437GAT(177)* 369GAT(113)* ; 488GAT(184)
g126 and 437GAT(177)* 369GAT(113)* ; 489GAT(185)
g127 and 437GAT(177)* 369GAT(113)* ; 490GAT(186)
g128 and 437GAT(177)* 369GAT(113)* ; 491GAT(187)
g129 and 432GAT(181) 310GAT(60) ; 476GAT(188)
g130 and 432GAT(181) 310GAT(60) ; 478GAT(189)
g131 and 432GAT(181) 310GAT(60) ; 480GAT(190)
g132 and 432GAT(181) 310GAT(60) ; 482GAT(191)
g133 and 445GAT(169)* 416GAT(144)* ; 495GAT(192)
g134 and 444GAT(170)* 413GAT(147)* ; 492GAT(193)
g135 and 427GAT(178) 153GAT(38) ; 481GAT(194)
g136 and 427GAT(178) 149GAT(36) ; 479GAT(195)
g137 and 427GAT(178) 146GAT(35) ; 477GAT(196)
g138 and 427GAT(178) 143GAT(34) ; 475GAT(197)
g139 and 426GAT(171)* 409GAT(150)* ; 463GAT(198)
g140 and 425GAT(172)* 406GAT(153)* ; 460GAT(199)
g141 and 424GAT(174) ; 451GAT(200)
g142 and 410GAT(160) 442GAT(175) ; 466GAT(201)
g143 and 1GAT(0) 443GAT(180) ; 483GAT(202)
g144 and 476GAT(188)* 475GAT(197)* ; 503GAT(203)
g145 and 478GAT(189)* 477GAT(196)* ; 505GAT(204)
g146 and 480GAT(190)* 479GAT(195)* ; 507GAT(205)
g147 and 482GAT(191)* 481GAT(194)* ; 509GAT(206)
g148 and 207GAT(48)* 495GAT(192)* ; 521GAT(207)
g149 and 207GAT(48) 495GAT(192) ; 520GAT(208)
g150 and 201GAT(47) 451GAT(200) ; 529GAT(209)
g151 and 195GAT(46) 451GAT(200) ; 528GAT(210)
g152 and 189GAT(45) 451GAT(200) ; 527GAT(211)
g153 and 183GAT(44) 451GAT(200) ; 526GAT(212)
g154 and 177GAT(43) 451GAT(200) ; 525GAT(213)
g155 and 171GAT(42) 451GAT(200) ; 524GAT(214)
g156 and 165GAT(41) 451GAT(200) ; 523GAT(215)
g157 and 159GAT(40) 451GAT(200) ; 522GAT(216)
g158 and 483GAT(202) 153GAT(38) ; 516GAT(217)
g159 and 483GAT(202) 149GAT(36) ; 514GAT(218)
g160 and 483GAT(202) 146GAT(35) ; 512GAT(219)
g161 and 483GAT(202) 143GAT(34) ; 510GAT(220)
g162 and 135GAT(32)* 463GAT(198)* ; 501GAT(221)
g163 and 135GAT(32) 463GAT(198) ; 500GAT(222)
g164 and 492GAT(193)* 130GAT(31)* ; 519GAT(223)
g165 and 492GAT(193) 130GAT(31) ; 518GAT(224)
g166 and 460GAT(199)* 130GAT(31)* ; 499GAT(225)
g167 and 460GAT(199) 130GAT(31) ; 498GAT(226)
g168 and 466GAT(201) 126GAT(30) ; 517GAT(227)
g169 and 466GAT(201) 121GAT(29) ; 515GAT(228)
g170 and 466GAT(201) 116GAT(28) ; 513GAT(229)
g171 and 466GAT(201) 111GAT(27) ; 511GAT(230)
g172 and 466GAT(201) 106GAT(26) ; 508GAT(231)
g173 and 466GAT(201) 101GAT(25) ; 506GAT(232)
g174 and 466GAT(201) 96GAT(24) ; 504GAT(233)
g175 and 466GAT(201) 91GAT(23) ; 502GAT(234)
g176 and 521GAT(207) 520GAT(208) ; 547GAT(235)
g177 and 517GAT(227)* 516GAT(217)* ; 543GAT(236)
g178 and 515GAT(228)* 514GAT(218)* ; 542GAT(237)
g179 and 513GAT(229)* 512GAT(219)* ; 541GAT(238)
g180 and 511GAT(230)* 510GAT(220)* ; 540GAT(239)
g181 and 508GAT(231)* 318GAT(72)* ; 539GAT(240)
g182 and 501GAT(221) 500GAT(222) ; 533GAT(241)
g183 and 519GAT(223) 518GAT(224) ; 544GAT(242)
g184 and 499GAT(225) 498GAT(226) ; 530GAT(243)
g185 and 504GAT(233)* 316GAT(93)* ; 537GAT(244)
g186 and 506GAT(232)* 317GAT(106)* ; 538GAT(245)
g187 and 502GAT(234)* 309GAT(107)* ; 536GAT(246)
g188 and 540GAT(239) 488GAT(184) ; 569GAT(247)
g189 and 541GAT(238) 489GAT(185) ; 573GAT(248)
g190 and 542GAT(237) 490GAT(186) ; 577GAT(249)
g191 and 543GAT(236) 491GAT(187) ; 581GAT(250)
g192 and 503GAT(203) 536GAT(246) ; 553GAT(251)
g193 and 505GAT(204) 537GAT(244) ; 557GAT(252)
g194 and 507GAT(205) 538GAT(245) ; 561GAT(253)
g195 and 509GAT(206) 539GAT(240) ; 565GAT(254)
g196 and 547GAT(235) ; 586GAT(255)
g197 and 547GAT(235) 544GAT(242) ; 587GAT(256)
g198 and 533GAT(241) ; 551GAT(257)
g199 and 533GAT(241) 530GAT(243) ; 552GAT(258)
g200 and 544GAT(242) ; 585GAT(259)
g201 and 530GAT(243) ; 550GAT(260)
g202 and 581GAT(250) 246GAT(53) ; 659GAT(261)
g203 and 577GAT(249) 246GAT(53) ; 650GAT(262)
g204 and 573GAT(248) 246GAT(53) ; 640GAT(263)
g205 and 569GAT(247) 246GAT(53) ; 631GAT(264)
g206 and 565GAT(254) 246GAT(53) ; 624GAT(265)
g207 and 561GAT(253) 246GAT(53) ; 615GAT(266)
g208 and 557GAT(252) 246GAT(53) ; 605GAT(267)
g209 and 553GAT(251) 246GAT(53) ; 596GAT(268)
g210 and 586GAT(255) 585GAT(259) ; 589GAT(269)
g211 and 201GAT(47)* 581GAT(250)* ; 654GAT(270)
g212 and 201GAT(47) 581GAT(250) ; 651GAT(271)
g213 and 195GAT(46)* 577GAT(249)* ; 644GAT(272)
g214 and 195GAT(46) 577GAT(249) ; 641GAT(273)
g215 and 189GAT(45)* 573GAT(248)* ; 635GAT(274)
g216 and 189GAT(45) 573GAT(248) ; 632GAT(275)
g217 and 183GAT(44)* 569GAT(247)* ; 628GAT(276)
g218 and 183GAT(44) 569GAT(247) ; 625GAT(277)
g219 and 177GAT(43)* 565GAT(254)* ; 619GAT(278)
g220 and 177GAT(43) 565GAT(254) ; 616GAT(279)
g221 and 171GAT(42)* 561GAT(253)* ; 609GAT(280)
g222 and 171GAT(42) 561GAT(253) ; 606GAT(281)
g223 and 165GAT(41)* 557GAT(252)* ; 600GAT(282)
g224 and 165GAT(41) 557GAT(252) ; 597GAT(283)
g225 and 159GAT(40)* 553GAT(251)* ; 593GAT(284)
g226 and 159GAT(40) 553GAT(251) ; 590GAT(285)
g227 and 551GAT(257) 550GAT(260) ; 588GAT(286)
g228 and 261GAT(57) 654GAT(270) 644GAT(272) 635GAT(274) ; 734GAT(287)
g229 and 261GAT(57) 654GAT(270) 644GAT(272) ; 733GAT(288)
g230 and 261GAT(57) 654GAT(270) ; 732GAT(289)
g231 and 659GAT(261)* 341GAT(61)* ; 731GAT(290)
g232 and 650GAT(262)* 339GAT(62)* ; 721GAT(291)
g233 and 640GAT(263)* 337GAT(63)* ; 712GAT(292)
g234 and 589GAT(269)* 587GAT(256)* ; 661GAT(293)
g235 and 651GAT(271) 654GAT(270) ; 727GAT(294)
g236 and 651GAT(271) ; 722GAT(295)
g237 and 641GAT(273) 644GAT(272) ; 717GAT(296)
g238 and 641GAT(273) ; 713GAT(297)
g239 and 632GAT(275) 635GAT(274) ; 708GAT(298)
g240 and 632GAT(275) ; 705GAT(299)
g241 and 625GAT(277) 628GAT(276) ; 700GAT(300)
g242 and 625GAT(277) ; 697GAT(301)
g243 and 526GAT(212)* 631GAT(264)* ; 704GAT(302)
g244 and 616GAT(279) 619GAT(278) ; 692GAT(303)
g245 and 616GAT(279) ; 687GAT(304)
g246 and 525GAT(213)* 624GAT(265)* ; 696GAT(305)
g247 and 606GAT(281) 609GAT(280) ; 682GAT(306)
g248 and 606GAT(281) ; 678GAT(307)
g249 and 524GAT(214)* 615GAT(266)* ; 686GAT(308)
g250 and 597GAT(283) 600GAT(282) ; 673GAT(309)
g251 and 597GAT(283) ; 670GAT(310)
g252 and 523GAT(215)* 605GAT(267)* ; 677GAT(311)
g253 and 590GAT(285) 593GAT(284) ; 665GAT(312)
g254 and 590GAT(285) ; 662GAT(313)
g255 and 522GAT(216)* 596GAT(268)* ; 669GAT(314)
g256 and 588GAT(286)* 552GAT(258)* ; 660GAT(315)
g257 and 261GAT(57) 727GAT(294) ; 758GAT(316)
g258 and 261GAT(57)* 727GAT(294)* ; 757GAT(317)
g259 and 722GAT(295) 237GAT(52) ; 760GAT(318)
g260 and 713GAT(297) 237GAT(52) ; 755GAT(319)
g261 and 705GAT(299) 237GAT(52) ; 752GAT(320)
g262 and 697GAT(301) 237GAT(52) ; 749GAT(321)
g263 and 687GAT(304) 237GAT(52) ; 746GAT(322)
g264 and 678GAT(307) 237GAT(52) ; 743GAT(323)
g265 and 670GAT(310) 237GAT(52) ; 740GAT(324)
g266 and 662GAT(313) 237GAT(52) ; 737GAT(325)
g267 and 727GAT(294) 228GAT(51) ; 759GAT(326)
g268 and 717GAT(296) 228GAT(51) ; 754GAT(327)
g269 and 708GAT(298) 228GAT(51) ; 751GAT(328)
g270 and 700GAT(300) 228GAT(51) ; 748GAT(329)
g271 and 692GAT(303) 228GAT(51) ; 745GAT(330)
g272 and 682GAT(306) 228GAT(51) ; 742GAT(331)
g273 and 673GAT(309) 228GAT(51) ; 739GAT(332)
g274 and 665GAT(312) 228GAT(51) ; 736GAT(333)
g275 and 661GAT(293) ; 768GAT(334)
g276 and 722GAT(295) ; 756GAT(335)
g277 and 722GAT(295) 644GAT(272) ; 761GAT(336)
g278 and 722GAT(295) 644GAT(272) 635GAT(274) ; 763GAT(337)
g279 and 713GAT(297) ; 753GAT(338)
g280 and 713GAT(297) 635GAT(274) ; 762GAT(339)
g281 and 705GAT(299) ; 750GAT(340)
g282 and 697GAT(301) ; 747GAT(341)
g283 and 687GAT(304) ; 744GAT(342)
g284 and 687GAT(304) 609GAT(280) ; 764GAT(343)
g285 and 687GAT(304) 609GAT(280) 600GAT(282) ; 766GAT(344)
g286 and 678GAT(307) ; 741GAT(345)
g287 and 678GAT(307) 600GAT(282) ; 765GAT(346)
g288 and 670GAT(310) ; 738GAT(347)
g289 and 662GAT(313) ; 735GAT(348)
g290 and 660GAT(315) ; 767GAT(349)
g291 and 758GAT(316)* 757GAT(317)* ; 786GAT(350)
g292 and 734GAT(287) 763GAT(337) 762GAT(339) 750GAT(340) ; 773GAT(351)
g293 and 733GAT(288) 761GAT(336) 753GAT(338) ; 778GAT(352)
g294 and 732GAT(289) 756GAT(335) ; 782GAT(353)
g295 and 760GAT(318)* 759GAT(326)* ; 787GAT(354)
g296 and 755GAT(319)* 754GAT(327)* ; 785GAT(355)
g297 and 752GAT(320)* 751GAT(328)* ; 781GAT(356)
g298 and 749GAT(321)* 748GAT(329)* ; 777GAT(357)
g299 and 746GAT(322)* 745GAT(330)* ; 772GAT(358)
g300 and 743GAT(323)* 742GAT(331)* ; 771GAT(359)
g301 and 740GAT(324)* 739GAT(332)* ; 770GAT(360)
g302 and 737GAT(325)* 736GAT(333)* ; 769GAT(361)
g303 and 786GAT(350) 219GAT(50) ; 794GAT(362)
g304 and 782GAT(353)* 717GAT(296)* ; 792GAT(363)
g305 and 782GAT(353) 717GAT(296) ; 793GAT(364)
g306 and 778GAT(352)* 708GAT(298)* ; 790GAT(365)
g307 and 778GAT(352) 708GAT(298) ; 791GAT(366)
g308 and 773GAT(351)* 700GAT(300)* ; 788GAT(367)
g309 and 773GAT(351) 700GAT(300) ; 789GAT(368)
g310 and 773GAT(351) 628GAT(276) ; 795GAT(369)
g311 and 793GAT(364)* 792GAT(363)* ; 804GAT(370)
g312 and 791GAT(366)* 790GAT(365)* ; 803GAT(371)
g313 and 789GAT(368)* 788GAT(367)* ; 802GAT(372)
g314 and 747GAT(341) 795GAT(369) ; 796GAT(373)
g315 and 794GAT(362)* 340GAT(73)* ; 805GAT(374)
g316 and 804GAT(370) 219GAT(50) ; 810GAT(375)
g317 and 803GAT(371) 219GAT(50) ; 809GAT(376)
g318 and 802GAT(372) 219GAT(50) ; 808GAT(377)
g319 and 529GAT(209) 731GAT(290) 787GAT(354) 805GAT(374) ; 811GAT(378)
g320 and 796GAT(373)* 692GAT(303)* ; 806GAT(379)
g321 and 796GAT(373) 692GAT(303) ; 807GAT(380)
g322 and 796GAT(373) 619GAT(278) ; 812GAT(381)
g323 and 796GAT(373) 619GAT(278) 609GAT(280) ; 813GAT(382)
g324 and 796GAT(373) 619GAT(278) 609GAT(280) 600GAT(282) ; 814GAT(383)
g325 and 811GAT(378) ; 829GAT(384)
g326 and 807GAT(380)* 806GAT(379)* ; 825GAT(385)
g327 and 812GAT(381) 744GAT(342) ; 822GAT(386)
g328 and 813GAT(382) 764GAT(343) 741GAT(345) ; 819GAT(387)
g329 and 814GAT(383) 766GAT(344) 765GAT(346) 738GAT(347) ; 815GAT(388)
g330 and 810GAT(375)* 338GAT(76)* ; 828GAT(389)
g331 and 809GAT(376)* 336GAT(77)* ; 827GAT(390)
g332 and 808GAT(377)* 335GAT(80)* ; 826GAT(391)
g333 and 825GAT(385) 219GAT(50) ; 836GAT(392)
g334 and 829GAT(384) ; 840GAT(393)
g335 and 528GAT(210) 721GAT(291) 785GAT(355) 828GAT(389) ; 839GAT(394)
g336 and 527GAT(211) 712GAT(292) 781GAT(356) 827GAT(390) ; 838GAT(395)
g337 and 704GAT(302) 777GAT(357) 826GAT(391) ; 837GAT(396)
g338 and 822GAT(386)* 682GAT(306)* ; 834GAT(397)
g339 and 822GAT(386) 682GAT(306) ; 835GAT(398)
g340 and 819GAT(387)* 673GAT(309)* ; 832GAT(399)
g341 and 819GAT(387) 673GAT(309) ; 833GAT(400)
g342 and 815GAT(388)* 665GAT(312)* ; 830GAT(401)
g343 and 815GAT(388) 665GAT(312) ; 831GAT(402)
g344 and 593GAT(284) 815GAT(388) ; 841GAT(403)
g345 and 840GAT(393) ; 850GAT(404)
g346 and 839GAT(394) ; 848GAT(405)
g347 and 838GAT(395) ; 847GAT(406)
g348 and 837GAT(396) ; 846GAT(407)
g349 and 835GAT(398)* 834GAT(397)* ; 844GAT(408)
g350 and 833GAT(400)* 832GAT(399)* ; 843GAT(409)
g351 and 831GAT(402)* 830GAT(401)* ; 842GAT(410)
g352 and 841GAT(403) 735GAT(348) ; 849GAT(411)
g353 and 836GAT(392)* 334GAT(81)* ; 845GAT(412)
g354 and 844GAT(408) 219GAT(50) ; 853GAT(413)
g355 and 843GAT(409) 219GAT(50) ; 852GAT(414)
g356 and 842GAT(410) 219GAT(50) ; 851GAT(415)
g357 and 848GAT(405) ; 857GAT(416)
g358 and 847GAT(406) ; 856GAT(417)
g359 and 846GAT(407) ; 855GAT(418)
g360 and 696GAT(305) 772GAT(358) 845GAT(412) ; 854GAT(419)
g361 and 849GAT(411) ; 858GAT(420)
g362 and 851GAT(415)* 417GAT(142)* ; 859GAT(421)
g363 and 857GAT(416) ; 865GAT(422)
g364 and 856GAT(417) ; 864GAT(423)
g365 and 855GAT(418) ; 863GAT(424)
g366 and 854GAT(419) ; 862GAT(425)
g367 and 858GAT(420) ; 866GAT(426)
g368 and 853GAT(413)* 333GAT(84)* ; 861GAT(427)
g369 and 852GAT(414)* 332GAT(85)* ; 860GAT(428)
g370 and 862GAT(425) ; 870GAT(429)
g371 and 686GAT(308) 771GAT(359) 861GAT(427) ; 869GAT(430)
g372 and 677GAT(311) 770GAT(360) 860GAT(428) ; 868GAT(431)
g373 and 669GAT(314) 769GAT(361) 859GAT(421) ; 867GAT(432)
g374 and 870GAT(429) ; 874GAT(433)
g375 and 869GAT(430) ; 873GAT(434)
g376 and 868GAT(431) ; 872GAT(435)
g377 and 867GAT(432) ; 871GAT(436)
g378 and 873GAT(434) ; 877GAT(437)
g379 and 872GAT(435) ; 876GAT(438)
g380 and 871GAT(436) ; 875GAT(439)
g381 and 877GAT(437) ; 880GAT(440)
g382 and 876GAT(438) ; 879GAT(441)
g383 and 875GAT(439) ; 878GAT(442)
g384 not 195GAT(46) ; 195GAT(46)*
g385 not 201GAT(47) ; 201GAT(47)*
g386 not 183GAT(44) ; 183GAT(44)*
g387 not 189GAT(45) ; 189GAT(45)*
g388 not 171GAT(42) ; 171GAT(42)*
g389 not 177GAT(43) ; 177GAT(43)*
g390 not 159GAT(40) ; 159GAT(40)*
g391 not 165GAT(41) ; 165GAT(41)*
g392 not 121GAT(29) ; 121GAT(29)*
g393 not 126GAT(30) ; 126GAT(30)*
g394 not 111GAT(27) ; 111GAT(27)*
g395 not 116GAT(28) ; 116GAT(28)*
g396 not 101GAT(25) ; 101GAT(25)*
g397 not 106GAT(26) ; 106GAT(26)*
g398 not 91GAT(23) ; 91GAT(23)*
g399 not 96GAT(24) ; 96GAT(24)*
g400 not 87GAT(19) ; 87GAT(19)*
g401 not 88GAT(20) ; 88GAT(20)*
g402 not 17GAT(3) ; 17GAT(3)*
g403 not 42GAT(7) ; 42GAT(7)*
g404 not 280GAT(108) ; 280GAT(108)*
g405 not 286GAT(92) ; 286GAT(92)*
g406 not 284GAT(95) ; 284GAT(95)*
g407 not 285GAT(102) ; 285GAT(102)*
g408 not 270GAT(111) ; 270GAT(111)*
g409 not 273GAT(103) ; 273GAT(103)*
g410 not 322GAT(105) ; 322GAT(105)*
g411 not 323GAT(104) ; 323GAT(104)*
g412 not 343GAT(135) ; 343GAT(135)*
g413 not 369GAT(113) ; 369GAT(113)*
g414 not 437GAT(177) ; 437GAT(177)*
g415 not 416GAT(144) ; 416GAT(144)*
g416 not 445GAT(169) ; 445GAT(169)*
g417 not 413GAT(147) ; 413GAT(147)*
g418 not 444GAT(170) ; 444GAT(170)*
g419 not 409GAT(150) ; 409GAT(150)*
g420 not 426GAT(171) ; 426GAT(171)*
g421 not 406GAT(153) ; 406GAT(153)*
g422 not 425GAT(172) ; 425GAT(172)*
g423 not 475GAT(197) ; 475GAT(197)*
g424 not 476GAT(188) ; 476GAT(188)*
g425 not 477GAT(196) ; 477GAT(196)*
g426 not 478GAT(189) ; 478GAT(189)*
g427 not 479GAT(195) ; 479GAT(195)*
g428 not 480GAT(190) ; 480GAT(190)*
g429 not 481GAT(194) ; 481GAT(194)*
g430 not 482GAT(191) ; 482GAT(191)*
g431 not 495GAT(192) ; 495GAT(192)*
g432 not 207GAT(48) ; 207GAT(48)*
g433 not 463GAT(198) ; 463GAT(198)*
g434 not 135GAT(32) ; 135GAT(32)*
g435 not 130GAT(31) ; 130GAT(31)*
g436 not 492GAT(193) ; 492GAT(193)*
g437 not 460GAT(199) ; 460GAT(199)*
g438 not 516GAT(217) ; 516GAT(217)*
g439 not 517GAT(227) ; 517GAT(227)*
g440 not 514GAT(218) ; 514GAT(218)*
g441 not 515GAT(228) ; 515GAT(228)*
g442 not 512GAT(219) ; 512GAT(219)*
g443 not 513GAT(229) ; 513GAT(229)*
g444 not 510GAT(220) ; 510GAT(220)*
g445 not 511GAT(230) ; 511GAT(230)*
g446 not 318GAT(72) ; 318GAT(72)*
g447 not 508GAT(231) ; 508GAT(231)*
g448 not 316GAT(93) ; 316GAT(93)*
g449 not 504GAT(233) ; 504GAT(233)*
g450 not 317GAT(106) ; 317GAT(106)*
g451 not 506GAT(232) ; 506GAT(232)*
g452 not 309GAT(107) ; 309GAT(107)*
g453 not 502GAT(234) ; 502GAT(234)*
g454 not 581GAT(250) ; 581GAT(250)*
g455 not 577GAT(249) ; 577GAT(249)*
g456 not 573GAT(248) ; 573GAT(248)*
g457 not 569GAT(247) ; 569GAT(247)*
g458 not 565GAT(254) ; 565GAT(254)*
g459 not 561GAT(253) ; 561GAT(253)*
g460 not 557GAT(252) ; 557GAT(252)*
g461 not 553GAT(251) ; 553GAT(251)*
g462 not 341GAT(61) ; 341GAT(61)*
g463 not 659GAT(261) ; 659GAT(261)*
g464 not 339GAT(62) ; 339GAT(62)*
g465 not 650GAT(262) ; 650GAT(262)*
g466 not 337GAT(63) ; 337GAT(63)*
g467 not 640GAT(263) ; 640GAT(263)*
g468 not 587GAT(256) ; 587GAT(256)*
g469 not 589GAT(269) ; 589GAT(269)*
g470 not 631GAT(264) ; 631GAT(264)*
g471 not 526GAT(212) ; 526GAT(212)*
g472 not 624GAT(265) ; 624GAT(265)*
g473 not 525GAT(213) ; 525GAT(213)*
g474 not 615GAT(266) ; 615GAT(266)*
g475 not 524GAT(214) ; 524GAT(214)*
g476 not 605GAT(267) ; 605GAT(267)*
g477 not 523GAT(215) ; 523GAT(215)*
g478 not 596GAT(268) ; 596GAT(268)*
g479 not 522GAT(216) ; 522GAT(216)*
g480 not 552GAT(258) ; 552GAT(258)*
g481 not 588GAT(286) ; 588GAT(286)*
g482 not 727GAT(294) ; 727GAT(294)*
g483 not 261GAT(57) ; 261GAT(57)*
g484 not 757GAT(317) ; 757GAT(317)*
g485 not 758GAT(316) ; 758GAT(316)*
g486 not 759GAT(326) ; 759GAT(326)*
g487 not 760GAT(318) ; 760GAT(318)*
g488 not 754GAT(327) ; 754GAT(327)*
g489 not 755GAT(319) ; 755GAT(319)*
g490 not 751GAT(328) ; 751GAT(328)*
g491 not 752GAT(320) ; 752GAT(320)*
g492 not 748GAT(329) ; 748GAT(329)*
g493 not 749GAT(321) ; 749GAT(321)*
g494 not 745GAT(330) ; 745GAT(330)*
g495 not 746GAT(322) ; 746GAT(322)*
g496 not 742GAT(331) ; 742GAT(331)*
g497 not 743GAT(323) ; 743GAT(323)*
g498 not 739GAT(332) ; 739GAT(332)*
g499 not 740GAT(324) ; 740GAT(324)*
g500 not 736GAT(333) ; 736GAT(333)*
g501 not 737GAT(325) ; 737GAT(325)*
g502 not 717GAT(296) ; 717GAT(296)*
g503 not 782GAT(353) ; 782GAT(353)*
g504 not 708GAT(298) ; 708GAT(298)*
g505 not 778GAT(352) ; 778GAT(352)*
g506 not 700GAT(300) ; 700GAT(300)*
g507 not 773GAT(351) ; 773GAT(351)*
g508 not 792GAT(363) ; 792GAT(363)*
g509 not 793GAT(364) ; 793GAT(364)*
g510 not 790GAT(365) ; 790GAT(365)*
g511 not 791GAT(366) ; 791GAT(366)*
g512 not 788GAT(367) ; 788GAT(367)*
g513 not 789GAT(368) ; 789GAT(368)*
g514 not 340GAT(73) ; 340GAT(73)*
g515 not 794GAT(362) ; 794GAT(362)*
g516 not 692GAT(303) ; 692GAT(303)*
g517 not 796GAT(373) ; 796GAT(373)*
g518 not 806GAT(379) ; 806GAT(379)*
g519 not 807GAT(380) ; 807GAT(380)*
g520 not 338GAT(76) ; 338GAT(76)*
g521 not 810GAT(375) ; 810GAT(375)*
g522 not 336GAT(77) ; 336GAT(77)*
g523 not 809GAT(376) ; 809GAT(376)*
g524 not 335GAT(80) ; 335GAT(80)*
g525 not 808GAT(377) ; 808GAT(377)*
g526 not 682GAT(306) ; 682GAT(306)*
g527 not 822GAT(386) ; 822GAT(386)*
g528 not 673GAT(309) ; 673GAT(309)*
g529 not 819GAT(387) ; 819GAT(387)*
g530 not 665GAT(312) ; 665GAT(312)*
g531 not 815GAT(388) ; 815GAT(388)*
g532 not 834GAT(397) ; 834GAT(397)*
g533 not 835GAT(398) ; 835GAT(398)*
g534 not 832GAT(399) ; 832GAT(399)*
g535 not 833GAT(400) ; 833GAT(400)*
g536 not 830GAT(401) ; 830GAT(401)*
g537 not 831GAT(402) ; 831GAT(402)*
g538 not 334GAT(81) ; 334GAT(81)*
g539 not 836GAT(392) ; 836GAT(392)*
g540 not 417GAT(142) ; 417GAT(142)*
g541 not 851GAT(415) ; 851GAT(415)*
g542 not 333GAT(84) ; 333GAT(84)*
g543 not 853GAT(413) ; 853GAT(413)*
g544 not 332GAT(85) ; 332GAT(85)*
g545 not 852GAT(414) ; 852GAT(414)*
