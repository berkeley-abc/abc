name C432.iscas
i 1GAT(0)
i 4GAT(1)
i 8GAT(2)
i 11GAT(3)
i 14GAT(4)
i 17GAT(5)
i 21GAT(6)
i 24GAT(7)
i 27GAT(8)
i 30GAT(9)
i 34GAT(10)
i 37GAT(11)
i 40GAT(12)
i 43GAT(13)
i 47GAT(14)
i 50GAT(15)
i 53GAT(16)
i 56GAT(17)
i 60GAT(18)
i 63GAT(19)
i 66GAT(20)
i 69GAT(21)
i 73GAT(22)
i 76GAT(23)
i 79GAT(24)
i 82GAT(25)
i 86GAT(26)
i 89GAT(27)
i 92GAT(28)
i 95GAT(29)
i 99GAT(30)
i 102GAT(31)
i 105GAT(32)
i 108GAT(33)
i 112GAT(34)
i 115GAT(35)

o 223GAT(84)
o 329GAT(133)
o 370GAT(163)
o 421GAT(188)
o 430GAT(193)
o 431GAT(194)
o 432GAT(195)

g1 and 108GAT(33) ; 151GAT(36)
g2 and 102GAT(31) ; 150GAT(37)
g3 and 95GAT(29) ; 147GAT(38)
g4 and 89GAT(27) ; 146GAT(39)
g5 and 82GAT(25) ; 143GAT(40)
g6 and 76GAT(23) ; 142GAT(41)
g7 and 69GAT(21) ; 139GAT(42)
g8 and 63GAT(19) ; 138GAT(43)
g9 and 56GAT(17) ; 135GAT(44)
g10 and 50GAT(15) ; 134GAT(45)
g11 and 43GAT(13) ; 131GAT(46)
g12 and 37GAT(11) ; 130GAT(47)
g13 and 30GAT(9) ; 127GAT(48)
g14 and 24GAT(7) ; 126GAT(49)
g15 and 17GAT(5) ; 123GAT(50)
g16 and 11GAT(3) ; 122GAT(51)
g17 and 4GAT(1) ; 119GAT(52)
g18 and 1GAT(0) ; 118GAT(53)
g19 and 151GAT(36)* 115GAT(35)* ; 198GAT(54)
g20 and 151GAT(36)* 112GAT(34)* ; 197GAT(55)
g21 and 108GAT(33) 150GAT(37) ; 180GAT(56)
g22 and 147GAT(38)* 105GAT(32)* ; 196GAT(57)
g23 and 147GAT(38)* 99GAT(30)* ; 195GAT(58)
g24 and 95GAT(29) 146GAT(39) ; 177GAT(59)
g25 and 143GAT(40)* 92GAT(28)* ; 194GAT(60)
g26 and 143GAT(40)* 86GAT(26)* ; 193GAT(61)
g27 and 82GAT(25) 142GAT(41) ; 174GAT(62)
g28 and 139GAT(42)* 79GAT(24)* ; 192GAT(63)
g29 and 139GAT(42)* 73GAT(22)* ; 191GAT(64)
g30 and 69GAT(21) 138GAT(43) ; 171GAT(65)
g31 and 135GAT(44)* 66GAT(20)* ; 190GAT(66)
g32 and 135GAT(44)* 60GAT(18)* ; 189GAT(67)
g33 and 56GAT(17) 134GAT(45) ; 168GAT(68)
g34 and 131GAT(46)* 53GAT(16)* ; 188GAT(69)
g35 and 131GAT(46)* 47GAT(14)* ; 187GAT(70)
g36 and 43GAT(13) 130GAT(47) ; 165GAT(71)
g37 and 127GAT(48)* 40GAT(12)* ; 186GAT(72)
g38 and 127GAT(48)* 34GAT(10)* ; 185GAT(73)
g39 and 30GAT(9) 126GAT(49) ; 162GAT(74)
g40 and 123GAT(50)* 27GAT(8)* ; 184GAT(75)
g41 and 123GAT(50)* 21GAT(6)* ; 183GAT(76)
g42 and 17GAT(5) 122GAT(51) ; 159GAT(77)
g43 and 119GAT(52)* 14GAT(4)* ; 158GAT(78)
g44 and 119GAT(52)* 8GAT(2)* ; 157GAT(79)
g45 and 4GAT(1) 118GAT(53) ; 154GAT(80)
g46 and 180GAT(56) 177GAT(59) 174GAT(62) 171GAT(65) 168GAT(68) 165GAT(71) 162GAT(74) 159GAT(77) 154GAT(80) ; 199GAT(81)
g47 and 199GAT(81) ; 203GAT(82)
g48 and 199GAT(81) ; 213GAT(83)
g49 and 199GAT(81) ; 223GAT(84)
g50 or internal__52 internal__51 ; 251GAT(85)
g51 and 180GAT(56) 203GAT(82)* ; internal__51
g52 and 180GAT(56)* 203GAT(82) ; internal__52
g53 and 102GAT(31) 213GAT(83) ; 259GAT(86)
g54 or internal__56 internal__55 ; 247GAT(87)
g55 and 177GAT(59) 203GAT(82)* ; internal__55
g56 and 177GAT(59)* 203GAT(82) ; internal__56
g57 and 89GAT(27) 213GAT(83) ; 258GAT(88)
g58 or internal__60 internal__59 ; 243GAT(89)
g59 and 174GAT(62) 203GAT(82)* ; internal__59
g60 and 174GAT(62)* 203GAT(82) ; internal__60
g61 and 76GAT(23) 213GAT(83) ; 257GAT(90)
g62 or internal__64 internal__63 ; 239GAT(91)
g63 and 171GAT(65) 203GAT(82)* ; internal__63
g64 and 171GAT(65)* 203GAT(82) ; internal__64
g65 and 63GAT(19) 213GAT(83) ; 256GAT(92)
g66 or internal__68 internal__67 ; 236GAT(93)
g67 and 168GAT(68) 203GAT(82)* ; internal__67
g68 and 168GAT(68)* 203GAT(82) ; internal__68
g69 and 50GAT(15) 213GAT(83) ; 255GAT(94)
g70 or internal__72 internal__71 ; 233GAT(95)
g71 and 165GAT(71) 203GAT(82)* ; internal__71
g72 and 165GAT(71)* 203GAT(82) ; internal__72
g73 and 37GAT(11) 213GAT(83) ; 254GAT(96)
g74 or internal__76 internal__75 ; 230GAT(97)
g75 and 162GAT(74) 203GAT(82)* ; internal__75
g76 and 162GAT(74)* 203GAT(82) ; internal__76
g77 and 24GAT(7) 213GAT(83) ; 250GAT(98)
g78 or internal__80 internal__79 ; 227GAT(99)
g79 and 159GAT(77) 203GAT(82)* ; internal__79
g80 and 159GAT(77)* 203GAT(82) ; internal__80
g81 and 11GAT(3) 213GAT(83) ; 246GAT(100)
g82 or internal__84 internal__83 ; 224GAT(101)
g83 and 154GAT(80) 203GAT(82)* ; internal__83
g84 and 154GAT(80)* 203GAT(82) ; internal__84
g85 and 213GAT(83) 1GAT(0) ; 242GAT(102)
g86 and 198GAT(54) 251GAT(85) ; 295GAT(103)
g87 and 197GAT(55) 251GAT(85) ; 285GAT(104)
g88 and 196GAT(57) 247GAT(87) ; 294GAT(105)
g89 and 195GAT(58) 247GAT(87) ; 282GAT(106)
g90 and 194GAT(60) 243GAT(89) ; 293GAT(107)
g91 and 193GAT(61) 243GAT(89) ; 279GAT(108)
g92 and 192GAT(63) 239GAT(91) ; 292GAT(109)
g93 and 191GAT(64) 239GAT(91) ; 276GAT(110)
g94 and 190GAT(66) 236GAT(93) ; 291GAT(111)
g95 and 189GAT(67) 236GAT(93) ; 273GAT(112)
g96 and 188GAT(69) 233GAT(95) ; 290GAT(113)
g97 and 187GAT(70) 233GAT(95) ; 270GAT(114)
g98 and 186GAT(72) 230GAT(97) ; 289GAT(115)
g99 and 185GAT(73) 230GAT(97) ; 267GAT(116)
g100 and 184GAT(75) 227GAT(99) ; 288GAT(117)
g101 and 183GAT(76) 227GAT(99) ; 264GAT(118)
g102 and 158GAT(78) 224GAT(101) ; 263GAT(119)
g103 and 157GAT(79) 224GAT(101) ; 260GAT(120)
g104 and 295GAT(103) ; 308GAT(121)
g105 and 285GAT(104) 282GAT(106) 279GAT(108) 276GAT(110) 273GAT(112) 270GAT(114) 267GAT(116) 264GAT(118) 260GAT(120) ; 296GAT(122)
g106 and 294GAT(105) ; 307GAT(123)
g107 and 293GAT(107) ; 306GAT(124)
g108 and 292GAT(109) ; 305GAT(125)
g109 and 291GAT(111) ; 304GAT(126)
g110 and 290GAT(113) ; 303GAT(127)
g111 and 289GAT(115) ; 302GAT(128)
g112 and 288GAT(117) ; 301GAT(129)
g113 and 263GAT(119) ; 300GAT(130)
g114 and 296GAT(122) ; 309GAT(131)
g115 and 296GAT(122) ; 319GAT(132)
g116 and 296GAT(122) ; 329GAT(133)
g117 and 112GAT(34) 319GAT(132) ; 347GAT(134)
g118 or internal__120 internal__119 ; 343GAT(135)
g119 and 285GAT(104) 309GAT(131)* ; internal__119
g120 and 285GAT(104)* 309GAT(131) ; internal__120
g121 and 99GAT(30) 319GAT(132) ; 346GAT(136)
g122 or internal__124 internal__123 ; 341GAT(137)
g123 and 282GAT(106) 309GAT(131)* ; internal__123
g124 and 282GAT(106)* 309GAT(131) ; internal__124
g125 and 86GAT(26) 319GAT(132) ; 345GAT(138)
g126 or internal__128 internal__127 ; 339GAT(139)
g127 and 279GAT(108) 309GAT(131)* ; internal__127
g128 and 279GAT(108)* 309GAT(131) ; internal__128
g129 and 73GAT(22) 319GAT(132) ; 344GAT(140)
g130 or internal__132 internal__131 ; 337GAT(141)
g131 and 276GAT(110) 309GAT(131)* ; internal__131
g132 and 276GAT(110)* 309GAT(131) ; internal__132
g133 and 60GAT(18) 319GAT(132) ; 342GAT(142)
g134 or internal__136 internal__135 ; 335GAT(143)
g135 and 273GAT(112) 309GAT(131)* ; internal__135
g136 and 273GAT(112)* 309GAT(131) ; internal__136
g137 and 47GAT(14) 319GAT(132) ; 340GAT(144)
g138 or internal__140 internal__139 ; 333GAT(145)
g139 and 270GAT(114) 309GAT(131)* ; internal__139
g140 and 270GAT(114)* 309GAT(131) ; internal__140
g141 and 34GAT(10) 319GAT(132) ; 338GAT(146)
g142 or internal__144 internal__143 ; 332GAT(147)
g143 and 267GAT(116) 309GAT(131)* ; internal__143
g144 and 267GAT(116)* 309GAT(131) ; internal__144
g145 and 21GAT(6) 319GAT(132) ; 336GAT(148)
g146 or internal__148 internal__147 ; 331GAT(149)
g147 and 264GAT(118) 309GAT(131)* ; internal__147
g148 and 264GAT(118)* 309GAT(131) ; internal__148
g149 and 319GAT(132) 8GAT(2) ; 334GAT(150)
g150 or internal__152 internal__151 ; 330GAT(151)
g151 and 260GAT(120) 309GAT(131)* ; internal__151
g152 and 260GAT(120)* 309GAT(131) ; internal__152
g153 and 308GAT(121) 343GAT(135) ; 356GAT(152)
g154 and 307GAT(123) 341GAT(137) ; 355GAT(153)
g155 and 306GAT(124) 339GAT(139) ; 354GAT(154)
g156 and 305GAT(125) 337GAT(141) ; 353GAT(155)
g157 and 304GAT(126) 335GAT(143) ; 352GAT(156)
g158 and 303GAT(127) 333GAT(145) ; 351GAT(157)
g159 and 302GAT(128) 332GAT(147) ; 350GAT(158)
g160 and 301GAT(129) 331GAT(149) ; 349GAT(159)
g161 and 300GAT(130) 330GAT(151) ; 348GAT(160)
g162 and 356GAT(152) 355GAT(153) 354GAT(154) 353GAT(155) 352GAT(156) 351GAT(157) 350GAT(158) 349GAT(159) 348GAT(160) ; 357GAT(161)
g163 and 357GAT(161) ; 360GAT(162)
g164 and 357GAT(161) ; 370GAT(163)
g165 and 115GAT(35) 360GAT(162) ; 379GAT(164)
g166 and 105GAT(32) 360GAT(162) ; 378GAT(165)
g167 and 92GAT(28) 360GAT(162) ; 377GAT(166)
g168 and 79GAT(24) 360GAT(162) ; 376GAT(167)
g169 and 66GAT(20) 360GAT(162) ; 375GAT(168)
g170 and 53GAT(16) 360GAT(162) ; 374GAT(169)
g171 and 40GAT(12) 360GAT(162) ; 373GAT(170)
g172 and 27GAT(8) 360GAT(162) ; 372GAT(171)
g173 and 360GAT(162) 14GAT(4) ; 371GAT(172)
g174 and 108GAT(33) 379GAT(164) 347GAT(134) 259GAT(86) ; 414GAT(173)
g175 and 95GAT(29) 378GAT(165) 346GAT(136) 258GAT(88) ; 411GAT(174)
g176 and 82GAT(25) 377GAT(166) 345GAT(138) 257GAT(90) ; 407GAT(175)
g177 and 69GAT(21) 376GAT(167) 344GAT(140) 256GAT(92) ; 404GAT(176)
g178 and 56GAT(17) 375GAT(168) 342GAT(142) 255GAT(94) ; 399GAT(177)
g179 and 43GAT(13) 374GAT(169) 340GAT(144) 254GAT(96) ; 393GAT(178)
g180 and 30GAT(9) 373GAT(170) 338GAT(146) 250GAT(98) ; 386GAT(179)
g181 and 17GAT(5) 372GAT(171) 336GAT(148) 246GAT(100) ; 381GAT(180)
g182 and 371GAT(172) 334GAT(150) 242GAT(102) 4GAT(1) ; 380GAT(181)
g183 and 414GAT(173) 411GAT(174) 407GAT(175) 404GAT(176) 399GAT(177) 393GAT(178) 386GAT(179) 381GAT(180) ; 416GAT(182)
g184 and 411GAT(174) ; 420GAT(183)
g185 and 407GAT(175) ; 419GAT(184)
g186 and 404GAT(176) ; 418GAT(185)
g187 and 393GAT(178) ; 417GAT(186)
g188 and 380GAT(181) ; 415GAT(187)
g189 and 416GAT(182)* 415GAT(187)* ; 421GAT(188)
g190 and 420GAT(183) 407GAT(175) 393GAT(178) 386GAT(179) ; 429GAT(189)
g191 and 399GAT(177) 418GAT(185) 393GAT(178) 386GAT(179) ; 425GAT(190)
g192 and 419GAT(184) 393GAT(178) 399GAT(177) ; 428GAT(191)
g193 and 417GAT(186) 386GAT(179) ; 422GAT(192)
g194 and 399GAT(177) 422GAT(192) 386GAT(179) 381GAT(180) ; 430GAT(193)
g195 and 428GAT(191) 425GAT(190) 386GAT(179) 381GAT(180) ; 431GAT(194)
g196 and 429GAT(189) 425GAT(190) 422GAT(192) 381GAT(180) ; 432GAT(195)
g197 not 115GAT(35) ; 115GAT(35)*
g198 not 151GAT(36) ; 151GAT(36)*
g199 not 112GAT(34) ; 112GAT(34)*
g200 not 105GAT(32) ; 105GAT(32)*
g201 not 147GAT(38) ; 147GAT(38)*
g202 not 99GAT(30) ; 99GAT(30)*
g203 not 92GAT(28) ; 92GAT(28)*
g204 not 143GAT(40) ; 143GAT(40)*
g205 not 86GAT(26) ; 86GAT(26)*
g206 not 79GAT(24) ; 79GAT(24)*
g207 not 139GAT(42) ; 139GAT(42)*
g208 not 73GAT(22) ; 73GAT(22)*
g209 not 66GAT(20) ; 66GAT(20)*
g210 not 135GAT(44) ; 135GAT(44)*
g211 not 60GAT(18) ; 60GAT(18)*
g212 not 53GAT(16) ; 53GAT(16)*
g213 not 131GAT(46) ; 131GAT(46)*
g214 not 47GAT(14) ; 47GAT(14)*
g215 not 40GAT(12) ; 40GAT(12)*
g216 not 127GAT(48) ; 127GAT(48)*
g217 not 34GAT(10) ; 34GAT(10)*
g218 not 27GAT(8) ; 27GAT(8)*
g219 not 123GAT(50) ; 123GAT(50)*
g220 not 21GAT(6) ; 21GAT(6)*
g221 not 14GAT(4) ; 14GAT(4)*
g222 not 119GAT(52) ; 119GAT(52)*
g223 not 8GAT(2) ; 8GAT(2)*
g224 not 203GAT(82) ; 203GAT(82)*
g225 not 180GAT(56) ; 180GAT(56)*
g226 not 177GAT(59) ; 177GAT(59)*
g227 not 174GAT(62) ; 174GAT(62)*
g228 not 171GAT(65) ; 171GAT(65)*
g229 not 168GAT(68) ; 168GAT(68)*
g230 not 165GAT(71) ; 165GAT(71)*
g231 not 162GAT(74) ; 162GAT(74)*
g232 not 159GAT(77) ; 159GAT(77)*
g233 not 154GAT(80) ; 154GAT(80)*
g234 not 309GAT(131) ; 309GAT(131)*
g235 not 285GAT(104) ; 285GAT(104)*
g236 not 282GAT(106) ; 282GAT(106)*
g237 not 279GAT(108) ; 279GAT(108)*
g238 not 276GAT(110) ; 276GAT(110)*
g239 not 273GAT(112) ; 273GAT(112)*
g240 not 270GAT(114) ; 270GAT(114)*
g241 not 267GAT(116) ; 267GAT(116)*
g242 not 264GAT(118) ; 264GAT(118)*
g243 not 260GAT(120) ; 260GAT(120)*
g244 not 415GAT(187) ; 415GAT(187)*
g245 not 416GAT(182) ; 416GAT(182)*
