name C5315.lsl
i 1P0
i 4P1
i 11P2
i 14P3
i 17P4
i 20P5
i 23P6
i 24P7
i 25P8
i 26P9
i 27P10
i 31P11
i 34P12
i 37P13
i 40P14
i 43P15
i 46P16
i 49P17
i 52P18
i 53P19
i 54P20
i 61P21
i 64P22
i 67P23
i 70P24
i 73P25
i 76P26
i 79P27
i 80P28
i 81P29
i 82P30
i 83P31
i 86P32
i 87P33
i 88P34
i 91P35
i 94P36
i 97P37
i 100P38
i 103P39
i 106P40
i 109P41
i 112P42
i 113P43
i 114P44
i 115P45
i 116P46
i 117P47
i 118P48
i 119P49
i 120P50
i 121P51
i 122P52
i 123P53
i 126P54
i 127P55
i 128P56
i 129P57
i 130P58
i 131P59
i 132P60
i 135P61
i 136P62
i 137P63
i 140P64
i 141P65
i 145P66
i 146P67
i 149P68
i 152P69
i 155P70
i 158P71
i 161P72
i 164P73
i 167P74
i 170P75
i 173P76
i 176P77
i 179P78
i 182P79
i 185P80
i 188P81
i 191P82
i 194P83
i 197P84
i 200P85
i 203P86
i 206P87
i 209P88
i 210P89
i 217P90
i 218P91
i 225P92
i 226P93
i 233P94
i 234P95
i 241P96
i 242P97
i 245P98
i 248P99
i 251P100
i 254P101
i 257P102
i 264P103
i 265P104
i 272P105
i 273P106
i 280P107
i 281P108
i 288P109
i 289P110
i 292P111
i 293P112
i 299P113
i 302P114
i 307P115
i 308P116
i 315P117
i 316P118
i 323P119
i 324P120
i 331P121
i 332P122
i 335P123
i 338P124
i 341P125
i 348P126
i 351P127
i 358P128
i 361P129
i 366P130
i 369P131
i 372P132
i 373P133
i 374P134
i 386P135
i 389P136
i 400P137
i 411P138
i 422P139
i 435P140
i 446P141
i 457P142
i 468P143
i 479P144
i 490P145
i 503P146
i 514P147
i 523P148
i 534P149
i 545P150
i 549P151
i 552P152
i 556P153
i 559P154
i 562P155
i 1497P156
i 1689P157
i 1690P158
i 1691P159
i 1694P160
i 2174P161
i 2358P162
i 2824P163
i 3173P164
i 3546P165
i 3548P166
i 3550P167
i 3552P168
i 3717P169
i 3724P170
i 4087P171
i 4088P172
i 4089P173
i 4090P174
i 4091P175
i 4092P176
i 4115P177
o 144P354
o 298P299
o 973P202
o 594P224
o 599P269
o 600P259
o 601P220
o 602P222
o 603P225
o 604P223
o 611P275
o 612P263
o 810P356
o 848P330
o 849P219
o 850P217
o 851P218
o 634P665
o 815P627
o 845P845
o 847P465
o 926P624
o 923P619
o 921P664
o 892P408
o 887P528
o 606P407
o 656P621
o 809P655
o 993P850
o 978P851
o 949P852
o 939P853
o 889P734
o 593P733
o 636P1280
o 704P1281
o 717P1282
o 820P1283
o 639P1275
o 673P1276
o 707P1277
o 715P1278
o 598P1623
o 610P1519
o 588P1696
o 615P1750
o 626P1752
o 632P1692
o 1002P1920
o 1004P1977
o 591P1894
o 618P1925
o 621P1893
o 629P1926
o 822P1933
o 838P2064
o 861P2070
o 623P2152
o 722P2131
o 832P2133
o 834P2123
o 836P2128
o 859P2132
o 871P2127
o 873P2124
o 875P2125
o 877P2126
o 998P2163
o 1000P2168
o 575P2240
o 585P2236
o 661P2178
o 693P2179
o 747P2187
o 752P2189
o 757P2190
o 762P2184
o 787P2186
o 792P2188
o 797P2191
o 802P2183
o 642P2222
o 664P2223
o 667P2224
o 670P2225
o 676P2229
o 696P2226
o 699P2227
o 702P2228
o 818P2273
o 813P2260
o 824P2274
o 826P2275
o 828P2233
o 830P2182
o 854P2268
o 863P2276
o 865P2277
o 867P2237
o 869P2181
o 712P2297
o 727P2298
o 732P2300
o 737P2279
o 742P2238
o 772P2299
o 777P2278
o 782P2239
o 645P2271
o 648P2295
o 651P2314
o 654P2315
o 679P2272
o 682P2296
o 685P2316
o 688P2317
o 843P2455
o 882P2456
o 767P2479
o 807P2480
o 658P2483
o 690P2484
g144P354 or 141P65 ; 144P354
g298P299 or 293P112 ; 298P299
g973P202 or 3173P164 ; 973P202
g594P224 or B3 ; 594P224
g599P269 or B4 ; 599P269
g600P259 or B5 ; 600P259
g601P220 or B6 ; 601P220
g602P222 or B7 ; 602P222
g603P225 or B8 ; 603P225
g604P223 or B9 ; 604P223
g611P275 or B10 ; 611P275
g612P263 or B11 ; 612P263
g810P356 or B12 ; 810P356
g848P330 or B13 ; 848P330
g849P219 or B14 ; 849P219
g850P217 or B15 ; 850P217
g851P218 or B16 ; 851P218
g634P665 or B17 ; 634P665
g815P627 or B18 ; 815P627
g845P845 or B19 ; 845P845
g847P465 or B20 ; 847P465
g926P624 or 137P63 ; 926P624
g923P619 or 141P65 ; 923P619
g921P664 or 1P0 ; 921P664
g892P408 or 549P151 ; 892P408
g887P528 or 299P113 ; 887P528
g606P407 or B26 ; 606P407
g656P621 or B27 ; 656P621
g809P655 or B28 ; 809P655
g993P850 or 1P0 ; 993P850
g978P851 or 1P0 ; 978P851
g949P852 or 1P0 ; 949P852
g939P853 or 1P0 ; 939P853
g889P734 or 299P113 ; 889P734
g593P733 or B34 ; 593P733
g636P1280 or B35 ; 636P1280
g704P1281 or B36 ; 704P1281
g717P1282 or B37 ; 717P1282
g820P1283 or B38 ; 820P1283
g639P1275 or B39 ; 639P1275
g673P1276 or B40 ; 673P1276
g707P1277 or B41 ; 707P1277
g715P1278 or B42 ; 715P1278
g598P1623 or B43 ; 598P1623
g610P1519 or B44 ; 610P1519
g588P1696 or B45 ; 588P1696
g615P1750 or B46 ; 615P1750
g626P1752 or B47 ; 626P1752
g632P1692 or B48 ; 632P1692
g1002P1920 or B49 ; 1002P1920
g1004P1977 or B50 ; 1004P1977
g591P1894 or B51 ; 591P1894
g618P1925 or B52 ; 618P1925
g621P1893 or B53 ; 621P1893
g629P1926 or B54 ; 629P1926
g822P1933 or B55 ; 822P1933
g838P2064 or B56 ; 838P2064
g861P2070 or B57 ; 861P2070
g623P2152 or B58 ; 623P2152
g722P2131 or B59 ; 722P2131
g832P2133 or B60 ; 832P2133
g834P2123 or B61 ; 834P2123
g836P2128 or B62 ; 836P2128
g859P2132 or B63 ; 859P2132
g871P2127 or B64 ; 871P2127
g873P2124 or B65 ; 873P2124
g875P2125 or B66 ; 875P2125
g877P2126 or B67 ; 877P2126
g998P2163 or B68 ; 998P2163
g1000P2168 or B69 ; 1000P2168
g575P2240 or B70 ; 575P2240
g585P2236 or B71 ; 585P2236
g661P2178 or B72 ; 661P2178
g693P2179 or B73 ; 693P2179
g747P2187 or B74 ; 747P2187
g752P2189 or B75 ; 752P2189
g757P2190 or B76 ; 757P2190
g762P2184 or B77 ; 762P2184
g787P2186 or B78 ; 787P2186
g792P2188 or B79 ; 792P2188
g797P2191 or B80 ; 797P2191
g802P2183 or B81 ; 802P2183
g642P2222 or B82 ; 642P2222
g664P2223 or B83 ; 664P2223
g667P2224 or B84 ; 667P2224
g670P2225 or B85 ; 670P2225
g676P2229 or B86 ; 676P2229
g696P2226 or B87 ; 696P2226
g699P2227 or B88 ; 699P2227
g702P2228 or B89 ; 702P2228
g818P2273 or B90 ; 818P2273
g813P2260 or B91 ; 813P2260
g824P2274 or B92 ; 824P2274
g826P2275 or B93 ; 826P2275
g828P2233 or B94 ; 828P2233
g830P2182 or B95 ; 830P2182
g854P2268 or B96 ; 854P2268
g863P2276 or B97 ; 863P2276
g865P2277 or B98 ; 865P2277
g867P2237 or B99 ; 867P2237
g869P2181 or B100 ; 869P2181
g712P2297 or B101 ; 712P2297
g727P2298 or B102 ; 727P2298
g732P2300 or B103 ; 732P2300
g737P2279 or B104 ; 737P2279
g742P2238 or B105 ; 742P2238
g772P2299 or B106 ; 772P2299
g777P2278 or B107 ; 777P2278
g782P2239 or B108 ; 782P2239
g645P2271 or B109 ; 645P2271
g648P2295 or B110 ; 648P2295
g651P2314 or B111 ; 651P2314
g654P2315 or B112 ; 654P2315
g679P2272 or B113 ; 679P2272
g682P2296 or B114 ; 682P2296
g685P2316 or B115 ; 685P2316
g688P2317 or B116 ; 688P2317
g843P2455 or B117 ; 843P2455
g882P2456 or B118 ; 882P2456
g767P2479 or B119 ; 767P2479
g807P2480 or B120 ; 807P2480
g658P2483 or B121 ; 658P2483
g690P2484 or B122 ; 690P2484
gB3 not 545P150 ; B3
gB4 not 348P126 ; B4
gB5 not 366P130 ; B5
gB6 and 552P152 562P155 ; B6
gB7 not 549P151 ; B7
gB8 not 545P150 ; B8
gB9 not 545P150 ; B9
gB10 not 338P124 ; B10
gB11 not 358P128 ; B11
gB12 and 141P65 145P66 ; B12
gB13 not 245P98 ; B13
gB14 not 552P152 ; B14
gB15 not 562P155 ; B15
gB16 not 559P154 ; B16
gB17 not 633P365 ; B17
g3173P164_b not 3173P164 ; 3173P164_b
gB18 and 136P62 3173P164_b ; B18
gB19 not 844P657 ; B19
gB20 not 846P254 ; B20
gB26 not 549P151 ; B26
g140P64_b not 140P64 ; 140P64_b
g2822P361_b not 2822P361 ; 2822P361_b
gB27 or 140P64_b 2822P361_b ; B27
gB28 not 2822P361 ; B28
gB34 not 299P113 ; B34
gB35 not 635P1114 ; B35
gB36 not 703P1115 ; B36
gB37 not 716P1116 ; B37
gB38 not 819P1117 ; B38
gB39 and 141P65 637P965 ; B39
gB40 and 141P65 671P966 ; B40
gB41 and 141P65 705P964 ; B41
gB42 and 141P65 713P967 ; B42
gB43 and 595P1463 596P1412 3328P916 ; B43
g3350P1331_b not 3350P1331 ; 3350P1331_b
gB44 and 607P1425 608P1440 3350P1331_b ; B44
gB45 and 1437P1530 1451P1551 ; B45
gB46 and 1843P1630 1857P1608 ; B46
gB47 and 2113P1632 2128P1619 ; B47
gB48 and 1166P1522 1179P1552 ; B48
g3532P1627_b not 3532P1627 ; 3532P1627_b
g3531P1757_b not 3531P1757 ; 3531P1757_b
gB49 or 3532P1627_b 3531P1757_b ; B49
g3967P1769_b not 3967P1769 ; 3967P1769_b
g3966P1862_b not 3966P1862 ; 3966P1862_b
gB50 or 3967P1769_b 3966P1862_b ; B50
gB51 or 589P1711 590P1806 ; B51
gB52 or 616P1763 617P1849 ; B52
gB53 or 619P1710 620P1800 ; B53
gB54 or 627P1764 628P1853 ; B54
gB55 not 3848P1864 ; B55
gB56 not 3849P2024 ; B56
gB57 not 3790P2025 ; B57
gB58 not 1936P2105 ; B58
gB59 or 718P1867 719P2030 720P848 721P646 ; B59
gB60 not 4082P2071 ; B60
gB61 not 3851P2063 ; B61
gB62 not 3850P2069 ; B62
gB63 or 855P1866 856P2029 857P849 858P647 ; B63
gB64 not 4024P2068 ; B64
gB65 not 3793P2065 ; B65
gB66 not 3792P2066 ; B66
gB67 not 3791P2067 ; B67
g3537P2019_b not 3537P2019 ; 3537P2019_b
g3536P2059_b not 3536P2059 ; 3536P2059_b
gB68 or 3537P2019_b 3536P2059_b ; B68
g3542P2023_b not 3542P2023 ; 3542P2023_b
g3541P2062_b not 3541P2062 ; 3541P2062_b
gB69 or 3542P2023_b 3541P2062_b ; B69
g1200P1934_b not 1200P1934 ; 1200P1934_b
g1238P1953_b not 1238P1953 ; 1238P1953_b
g1248P1959_b not 1248P1959 ; 1248P1959_b
g1253P1960_b not 1253P1960 ; 1253P1960_b
g1243P1961_b not 1243P1961 ; 1243P1961_b
g1273P2005_b not 1273P2005 ; 1273P2005_b
g1268P2050_b not 1268P2050 ; 1268P2050_b
g1263P2111_b not 1263P2111 ; 1263P2111_b
g1258P2112_b not 1258P2112 ; 1258P2112_b
gB70 and 1200P1934_b 1238P1953_b 1248P1959_b 1253P1960_b 1243P1961_b 1273P2005_b 1268P2050_b 1263P2111_b 1258P2112_b ; B70
g1936P2105_b not 1936P2105 ; 1936P2105_b
g1878P1647_b not 1878P1647 ; 1878P1647_b
g1931P1914_b not 1931P1914 ; 1931P1914_b
g1926P1937_b not 1926P1937 ; 1926P1937_b
g1921P1939_b not 1921P1939 ; 1921P1939_b
g1916P1940_b not 1916P1940 ; 1916P1940_b
g1954P1997_b not 1954P1997 ; 1954P1997_b
g1949P2040_b not 1949P2040 ; 1949P2040_b
g1944P2104_b not 1944P2104 ; 1944P2104_b
gB71 and 1936P2105_b 1878P1647_b 1931P1914_b 1926P1937_b 1921P1939_b 1916P1940_b 1954P1997_b 1949P2040_b 1944P2104_b ; B71
gB72 and 137P63 659P2121 ; B72
gB73 and 137P63 691P2122 ; B73
gB74 or 743P2082 744P2081 745P841 746P654 ; B74
gB75 or 748P2086 749P2083 750P831 751P659 ; B75
gB76 or 753P2087 754P2084 755P832 756P660 ; B76
gB77 or 758P2031 759P2085 760P835 761P643 ; B77
gB78 or 783P2074 784P2077 785P840 786P653 ; B78
gB79 or 788P2075 789P2078 790P830 791P658 ; B79
gB80 or 793P2076 794P2079 795P833 796P661 ; B80
gB81 or 798P2028 799P2080 800P834 801P642 ; B81
gB82 and 137P63 640P2170 ; B82
gB83 and 137P63 662P2173 ; B83
gB84 and 137P63 665P2174 ; B84
gB85 and 137P63 668P2177 ; B85
gB86 and 137P63 674P2171 ; B86
gB87 and 137P63 694P2172 ; B87
gB88 and 137P63 697P2175 ; B88
gB89 and 137P63 700P2176 ; B89
g4114P359_b not 4114P359 ; 4114P359_b
gB90 and 817P2230 4114P359_b ; B90
gB91 or 811P2219 812P2205 ; B91
gB92 not 4086P2231 ; B92
gB93 not 4085P2232 ; B93
gB94 not 4084P2180 ; B94
gB95 not 4083P2130 ; B95
gB96 and 245P98 852P255 853P2202 ; B96
gB97 not 4028P2234 ; B97
gB98 not 4027P2235 ; B98
gB99 not 4026P2185 ; B99
gB100 not 4025P2129 ; B100
gB101 or 708P2243 709P2245 710P822 711P630 ; B101
gB102 or 723P2249 724P2247 725P823 726P631 ; B102
gB103 or 728P2250 729P2248 730P839 731P650 ; B103
gB104 or 733P2197 734P2196 735P825 736P633 ; B104
gB105 or 738P2141 739P2140 740P827 741P651 ; B105
gB106 or 768P2244 769P2246 770P838 771P649 ; B106
gB107 or 773P2194 774P2195 775P824 776P632 ; B107
gB108 or 778P2138 779P2139 780P826 781P652 ; B108
gB109 and 137P63 643P2221 ; B109
gB110 and 137P63 646P2269 ; B110
gB111 and 137P63 649P2292 ; B111
gB112 and 137P63 652P2293 ; B112
gB113 and 137P63 677P2220 ; B113
gB114 and 137P63 680P2270 ; B114
gB115 and 137P63 683P2291 ; B115
gB116 and 137P63 686P2294 ; B116
gB117 or 839P2241 840P2451 841P813 842P368 ; B117
gB118 or 878P2242 879P2452 880P815 881P370 ; B118
gB119 or 763P2472 764P2471 765P847 766P644 ; B119
gB120 or 803P2469 804P2470 805P846 806P645 ; B120
gB121 not 657P2481 ; B121
gB122 not 689P2482 ; B122
g1P0_b not 1P0 ; 1P0_b
g373P133_b not 373P133 ; 373P133_b
g633P365 or 1P0_b 373P133_b ; 633P365
g2824P163_b not 2824P163 ; 2824P163_b
g844P657 and 27P10 2824P163_b ; 844P657
g846P254 and 386P135 556P153 ; 846P254
g2822P361 and 27P10 31P11 ; 2822P361
g635P1114 and 3176P362 3197P953 ; 635P1114
g703P1115 and 3176P362 3200P952 ; 703P1115
g716P1116 and 3176P362 3203P951 ; 716P1116
g819P1117 and 3176P362 3194P954 ; 819P1117
g637P965 or 2881P678 2880P684 2879P960 2878P961 ; 637P965
g671P966 or 2877P679 2876P683 2875P956 2874P959 ; 671P966
g705P964 or 2869P677 2868P681 2866P958 2867P962 ; 705P964
g713P967 or 2873P680 2872P682 2870P955 2871P957 ; 713P967
g2933P933_b not 2933P933 ; 2933P933_b
g2942P1137_b not 2942P1137 ; 2942P1137_b
g2939P1144_b not 2939P1144 ; 2939P1144_b
g595P1463 and 2908P930 2933P933_b 2942P1137_b 2939P1144_b ; 595P1463
g3015P863_b not 3015P863 ; 3015P863_b
g3021P1123_b not 3021P1123 ; 3021P1123_b
g3018P1126_b not 3018P1126 ; 3018P1126_b
g3012P1132_b not 3012P1132 ; 3012P1132_b
g596P1412 and 3015P863_b 3021P1123_b 3018P1126_b 3012P1132_b ; 596P1412
g2615P1155_b not 2615P1155 ; 2615P1155_b
g2611P1159_b not 2611P1159 ; 2611P1159_b
g2623P1167_b not 2623P1167 ; 2623P1167_b
g2619P1171_b not 2619P1171 ; 2619P1171_b
g607P1425 and 2615P1155_b 2611P1159_b 2623P1167_b 2619P1171_b ; 607P1425
g2713P1178_b not 2713P1178 ; 2713P1178_b
g2709P1183_b not 2709P1183 ; 2709P1183_b
g2705P1186_b not 2705P1186 ; 2705P1186_b
g2717P1191_b not 2717P1191 ; 2717P1191_b
g608P1440 and 2713P1178_b 2709P1183_b 2705P1186_b 2717P1191_b ; 608P1440
g1437P1530 and 1307P1427 1289P1428 1278P1433 1422P1439 ; 1437P1530
g1451P1551 and 1332P1435 1390P1443 1365P1445 1344P1449 1430P1451 ; 1451P1551
g3165P927_b not 3165P927 ; 3165P927_b
g3167P931_b not 3167P931 ; 3167P931_b
g1843P1630 and 3165P927_b 3167P931_b 1758P1420 1730P1422 ; 1843P1630
g3137P914_b not 3137P914 ; 3137P914_b
g1857P1608 and 3137P914_b 1778P1307 1812P1404 1794P1406 1767P1417 ; 1857P1608
g2113P1632 and 3165P927_b 3167P931_b 2099P1419 1984P1423 ; 2113P1632
g2128P1619 and 3137P914_b 2021P1306 2067P1403 2042P1408 2009P1416 ; 2128P1619
g1166P1522 and 1052P1426 1034P1429 1023P1432 1080P1438 ; 1166P1522
g1179P1552 and 1089P1436 1134P1442 1116P1446 1100P1448 1152P1452 ; 1179P1552
g589P1711 or 1286P1007 1440P1534 1439P1539 1441P1563 ; 589P1711
g590P1806 and 1437P1530 1458P1719 ; 590P1806
g616P1763 or 3167P931 1846P1147 1845P1226 1847P1509 ; 616P1763
g617P1849 and 1843P1630 1863P1675 ; 617P1849
g619P1710 or 1031P1006 1169P1525 1168P1542 1170P1555 ; 619P1710
g620P1800 and 1166P1522 1185P1721 ; 620P1800
g627P1764 or 3167P931 2116P1152 2115P1229 2117P1504 ; 627P1764
g628P1853 and 2113P1632 2135P1673 ; 628P1853
g3848P1864 or 3838P804 3836P1120 3837P1653 ; 3848P1864
g3849P2024 or 3841P806 3839P1291 3840P1935 ; 3849P2024
g3790P2025 or 3780P816 3778P1293 3779P1936 ; 3790P2025
g1936P2105 or 1935P1994 1934P2039 ; 1936P2105
g4087P171_b not 4087P171 ; 4087P171_b
g4088P172_b not 4088P172 ; 4088P172_b
g718P1867 and 4087P171_b 4088P172_b 3848P1864 ; 718P1867
g719P2030 and 4087P171_b 4088P172 3790P2025 ; 719P2030
g720P848 and 11P2 4087P171 4088P172_b ; 720P848
g721P646 and 61P21 4087P171 4088P172 ; 721P646
g4082P2071 or 4069P837 4067P1284 4068P1980 ; 4082P2071
g3851P2063 or 3847P805 3845P963 3846P1982 ; 3851P2063
g3850P2069 or 3844P814 3842P1292 3843P1983 ; 3850P2069
g4089P173_b not 4089P173 ; 4089P173_b
g4090P174_b not 4090P174 ; 4090P174_b
g855P1866 and 4089P173_b 4090P174_b 3848P1864 ; 855P1866
g856P2029 and 4089P173 4090P174_b 3790P2025 ; 856P2029
g857P849 and 11P2 4089P173_b 4090P174 ; 857P849
g858P647 and 61P21 4089P173 4090P174 ; 858P647
g4024P2068 or 4011P811 4009P1287 4010P1981 ; 4024P2068
g3793P2065 or 3789P807 3787P1296 3788P1984 ; 3793P2065
g3792P2066 or 3786P808 3784P1295 3785P1985 ; 3792P2066
g3791P2067 or 3783P809 3781P1294 3782P1986 ; 3791P2067
g659P2121 or 1668P599 1667P797 1664P1870 1666P2035 ; 659P2121
g691P2122 or 2339P600 2338P796 2335P1869 2337P2033 ; 691P2122
g743P2082 and 4087P171_b 4088P172_b 4082P2071 ; 743P2082
g744P2081 and 4087P171_b 4088P172 4024P2068 ; 744P2081
g745P841 and 43P15 4087P171 4088P172_b ; 745P841
g746P654 and 37P13 4087P171 4088P172 ; 746P654
g748P2086 and 4087P171_b 4088P172_b 3851P2063 ; 748P2086
g749P2083 and 4087P171_b 4088P172 3793P2065 ; 749P2083
g750P831 and 76P26 4087P171 4088P172_b ; 750P831
g751P659 and 20P5 4087P171 4088P172 ; 751P659
g753P2087 and 4087P171_b 4088P172_b 3850P2069 ; 753P2087
g754P2084 and 4087P171_b 4088P172 3792P2066 ; 754P2084
g755P832 and 73P25 4087P171 4088P172_b ; 755P832
g756P660 and 17P4 4087P171 4088P172 ; 756P660
g758P2031 and 4087P171_b 4088P172_b 3849P2024 ; 758P2031
g759P2085 and 4087P171_b 4088P172 3791P2067 ; 759P2085
g760P835 and 67P23 4087P171 4088P172_b ; 760P835
g761P643 and 70P24 4087P171 4088P172 ; 761P643
g783P2074 and 4089P173_b 4090P174_b 4082P2071 ; 783P2074
g784P2077 and 4089P173 4090P174_b 4024P2068 ; 784P2077
g785P840 and 43P15 4089P173_b 4090P174 ; 785P840
g786P653 and 37P13 4089P173 4090P174 ; 786P653
g788P2075 and 4089P173_b 4090P174_b 3851P2063 ; 788P2075
g789P2078 and 4089P173 4090P174_b 3793P2065 ; 789P2078
g790P830 and 76P26 4089P173_b 4090P174 ; 790P830
g791P658 and 20P5 4089P173 4090P174 ; 791P658
g793P2076 and 4089P173_b 4090P174_b 3850P2069 ; 793P2076
g794P2079 and 4089P173 4090P174_b 3792P2066 ; 794P2079
g795P833 and 73P25 4089P173_b 4090P174 ; 795P833
g796P661 and 17P4 4089P173 4090P174 ; 796P661
g798P2028 and 4089P173_b 4090P174_b 3849P2024 ; 798P2028
g799P2080 and 4089P173 4090P174_b 3791P2067 ; 799P2080
g800P834 and 67P23 4089P173_b 4090P174 ; 800P834
g801P642 and 70P24 4089P173 4090P174 ; 801P642
g640P2170 or 1580P605 1579P787 1576P2097 1578P2101 ; 640P2170
g662P2173 or 1674P614 1673P794 1670P2034 1672P2100 ; 662P2173
g665P2174 or 1680P615 1679P801 1676P2095 1678P2099 ; 665P2174
g668P2177 or 1686P618 1685P802 1682P2096 1684P2098 ; 668P2177
g674P2171 or 2254P606 2253P786 2250P2090 2252P2094 ; 674P2171
g694P2172 or 2345P613 2344P795 2341P2032 2343P2093 ; 694P2172
g697P2175 or 2351P616 2350P800 2347P2088 2349P2092 ; 697P2175
g700P2176 or 2357P617 2356P803 2353P2089 2355P2091 ; 700P2176
g817P2230 or 3734P629 3731P1121 3733P1868 3735P2142 ; 817P2230
g811P2219 and 4113P1859 4096P2167 ; 811P2219
g812P2205 and 1936P2105 4096P2167 ; 812P2205
g4086P2231 or 4081P810 4079P1119 4080P2134 ; 4086P2231
g4085P2232 or 4078P812 4076P1118 4077P2135 ; 4085P2232
g4084P2180 or 4075P817 4073P1286 4074P2072 ; 4084P2180
g4083P2130 or 4072P821 4070P1285 4071P2026 ; 4083P2130
g852P255 and 386P135 552P152 556P153 559P154 ; 852P255
gB49_b not B49 ; B49_b
gB50_b not B50 ; B50_b
gB68_b not B68 ; B68_b
gB69_b not B69 ; B69_b
g853P2202 and 562P155 B49_b B50_b B68_b B69_b ; 853P2202
g4028P2234 or 4023P818 4021P1401 4022P2136 ; 4028P2234
g4027P2235 or 4020P819 4018P1290 4019P2137 ; 4027P2235
g4026P2185 or 4017P836 4015P1289 4016P2073 ; 4026P2185
g4025P2129 or 4014P820 4012P1288 4013P2027 ; 4025P2129
g708P2243 and 4089P173_b 4090P174_b 4086P2231 ; 708P2243
g709P2245 and 4089P173 4090P174_b 4028P2234 ; 709P2245
g710P822 and 109P41 4089P173_b 4090P174 ; 710P822
g711P630 and 106P40 4089P173 4090P174 ; 711P630
g723P2249 and 4087P171_b 4088P172_b 4086P2231 ; 723P2249
g724P2247 and 4087P171_b 4088P172 4028P2234 ; 724P2247
g725P823 and 109P41 4087P171 4088P172_b ; 725P823
g726P631 and 106P40 4087P171 4088P172 ; 726P631
g728P2250 and 4087P171_b 4088P172_b 4085P2232 ; 728P2250
g729P2248 and 4087P171_b 4088P172 4027P2235 ; 729P2248
g730P839 and 46P16 4087P171 4088P172_b ; 730P839
g731P650 and 49P17 4087P171 4088P172 ; 731P650
g733P2197 and 4087P171_b 4088P172_b 4084P2180 ; 733P2197
g734P2196 and 4087P171_b 4088P172 4026P2185 ; 734P2196
g735P825 and 100P38 4087P171 4088P172_b ; 735P825
g736P633 and 103P39 4087P171 4088P172 ; 736P633
g738P2141 and 4087P171_b 4088P172_b 4083P2130 ; 738P2141
g739P2140 and 4087P171_b 4088P172 4025P2129 ; 739P2140
g740P827 and 91P35 4087P171 4088P172_b ; 740P827
g741P651 and 40P14 4087P171 4088P172 ; 741P651
g768P2244 and 4089P173_b 4090P174_b 4085P2232 ; 768P2244
g769P2246 and 4089P173 4090P174_b 4027P2235 ; 769P2246
g770P838 and 46P16 4089P173_b 4090P174 ; 770P838
g771P649 and 49P17 4089P173 4090P174 ; 771P649
g773P2194 and 4089P173_b 4090P174_b 4084P2180 ; 773P2194
g774P2195 and 4089P173 4090P174_b 4026P2185 ; 774P2195
g775P824 and 100P38 4089P173_b 4090P174 ; 775P824
g776P632 and 103P39 4089P173 4090P174 ; 776P632
g778P2138 and 4089P173_b 4090P174_b 4083P2130 ; 778P2138
g779P2139 and 4089P173 4090P174_b 4025P2129 ; 779P2139
g780P826 and 91P35 4089P173_b 4090P174 ; 780P826
g781P652 and 40P14 4089P173 4090P174 ; 781P652
g643P2221 or 1586P604 1585P785 1582P2145 1584P2146 ; 643P2221
g646P2269 or 1592P607 1591P789 1588P2200 1590P2201 ; 646P2269
g649P2292 or 1598P610 1597P791 1594P2255 1596P2258 ; 649P2292
g652P2293 or 1604P611 1603P793 1600P2256 1602P2257 ; 652P2293
g677P2220 or 2260P603 2259P784 2256P2143 2258P2144 ; 677P2220
g680P2270 or 2266P608 2265P788 2262P2198 2264P2199 ; 680P2270
g683P2291 or 2272P609 2271P790 2268P2251 2270P2254 ; 683P2291
g686P2294 or 2278P612 2277P792 2274P2252 2276P2253 ; 686P2294
g4091P175_b not 4091P175 ; 4091P175_b
g4092P176_b not 4092P176 ; 4092P176_b
g3965P2153_b not 3965P2153 ; 3965P2153_b
g839P2241 and 4091P175_b 4092P176_b 3965P2153_b ; 839P2241
g840P2451 and 4091P175 4092P176_b 2198P2449 ; 840P2451
g841P813 and 120P50 4091P175_b 4092P176 ; 841P813
g842P368 and 4091P175 4092P176 ; 842P368
g3962P2154_b not 3962P2154 ; 3962P2154_b
g878P2242 and 4091P175_b 4092P176_b 3962P2154_b ; 878P2242
g879P2452 and 4091P175 4092P176_b 1521P2450 ; 879P2452
g880P815 and 118P48 4091P175_b 4092P176 ; 880P815
g881P370 and 4091P175 4092P176 ; 881P370
g763P2472 and 4087P171_b 4088P172_b 3656P2467 ; 763P2472
g764P2471 and 4087P171_b 4088P172 3655P2465 ; 764P2471
g765P847 and 14P3 4087P171 4088P172_b ; 765P847
g766P644 and 64P22 4087P171 4088P172 ; 766P644
g803P2469 and 4089P173_b 4090P174_b 3656P2467 ; 803P2469
g804P2470 and 4089P173 4090P174_b 3655P2465 ; 804P2470
g805P846 and 14P3 4089P173_b 4090P174 ; 805P846
g806P645 and 64P22 4089P173 4090P174 ; 806P645
g657P2481 and 137P63 1662P2477 ; 657P2481
g689P2482 and 137P63 2333P2478 ; 689P2482
g4114P359 and 135P61 4115P177 ; 4114P359
g3176P362 and 27P10 31P11 ; 3176P362
g3546P165_b not 3546P165 ; 3546P165_b
g2590P386 and 210P89 3546P165_b ; 2590P386
g2595P387 and 218P91 3546P165_b ; 2595P387
g2600P388 and 226P93 3546P165_b ; 2600P388
g2605P389 and 234P95 3546P165_b ; 2605P389
g2684P390 and 257P102 3546P165_b ; 2684P390
g2689P391 and 265P104 3546P165_b ; 2689P391
g2694P392 and 273P106 3546P165_b ; 2694P392
g2699P393 and 281P108 3546P165_b ; 2699P393
g2994P394 and 324P120 3546P165_b ; 2994P394
g3001P395 and 341P125 3546P165_b ; 3001P395
g3006P396 and 351P127 3546P165_b ; 3006P396
g3238P409 and 248P99 351P127 534P149 ; 3238P409
g3552P168_b not 3552P168 ; 3552P168_b
g2988P410 and 351P127 534P149 3552P168_b ; 2988P410
g2982P413 and 341P125 523P148 3552P168_b ; 2982P413
g3234P414 and 248P99 341P125 523P148 ; 3234P414
g3247P417 or 242P97 514P147 ; 3247P417
g3232P418 and 248P99 514P147 ; 3232P418
g2999P419 or 514P147 3546P165_b ; 2999P419
g2979P420 and 514P147 3552P168_b ; 2979P420
g2973P423 and 324P120 503P146 3552P168_b ; 2973P423
g3228P424 and 248P99 324P120 503P146 ; 3228P424
g3287P427 and 248P99 316P118 490P145 ; 3287P427
g2913P428 and 248P99 316P118 490P145 ; 2913P428
g2909P431 and 248P99 308P116 479P144 ; 2909P431
g3283P432 and 248P99 308P116 479P144 ; 3283P432
g3390P435 and 218P91 248P99 468P143 ; 3390P435
g2572P436 and 218P91 468P143 3552P168_b ; 2572P436
g3386P439 and 210P89 248P99 457P142 ; 3386P439
g2566P440 and 210P89 457P142 3552P168_b ; 2566P440
g3398P445 and 234P95 248P99 435P140 ; 3398P445
g2584P446 and 234P95 435P140 3552P168_b ; 2584P446
g3394P449 and 226P93 248P99 422P139 ; 3394P449
g2578P450 and 226P93 422P139 3552P168_b ; 2578P450
g2672P453 and 273P106 411P138 3552P168_b ; 2672P453
g3064P454 and 248P99 273P106 411P138 ; 3064P454
g3060P457 and 248P99 265P104 400P137 ; 3060P457
g2666P458 and 265P104 400P137 3552P168_b ; 2666P458
g2660P461 and 257P102 389P136 3552P168_b ; 2660P461
g3056P462 and 248P99 257P102 389P136 ; 3056P462
g3068P466 and 248P99 281P108 374P134 ; 3068P466
g2678P467 and 281P108 374P134 3552P168_b ; 2678P467
g3119P470 and 332P122 372P132 ; 3119P470
g3121P472 and 332P122 366P130 ; 3121P472
g3333P473 and 248P99 361P129 ; 3333P473
g3326P475 and 248P99 361P129 ; 3326P475
g3123P478 and 332P122 358P128 ; 3123P478
g3253P480 and 242P97 351P127 ; 3253P480
g3125P485 and 332P122 348P126 ; 3125P485
g3249P486 and 242P97 341P125 ; 3249P486
g3126P492 and 332P122 338P124 ; 3126P492
g3128P497 and 331P121 332P122 ; 3128P497
g3243P498 and 242P97 324P120 ; 3243P498
g3130P505 and 323P119 332P122 ; 3130P505
g3299P507 and 242P97 316P118 ; 3299P507
g2927P510 and 242P97 316P118 ; 2927P510
g3132P513 and 315P117 332P122 ; 3132P513
g3295P515 and 242P97 308P116 ; 3295P515
g2922P518 and 242P97 308P116 ; 2922P518
g3134P521 and 307P115 332P122 ; 3134P521
g3280P522 and 248P99 302P114 ; 3280P522
g2906P525 and 248P99 302P114 ; 2906P525
g3136P529 and 299P113 332P122 ; 3136P529
g3292P531 and 242P97 293P112 ; 3292P531
g2918P533 and 242P97 293P112 ; 2918P533
g2748P535 and 292P111 335P123 ; 2748P535
g2750P537 and 288P109 335P123 ; 2750P537
g3088P539 and 242P97 281P108 ; 3088P539
g2752P544 and 280P107 335P123 ; 2752P544
g3083P545 and 242P97 273P106 ; 3083P545
g2754P551 and 272P105 335P123 ; 2754P551
g3078P553 and 242P97 265P104 ; 3078P553
g2756P558 and 264P103 335P123 ; 2756P558
g3073P560 and 242P97 257P102 ; 3073P560
g3403P565 and 210P89 242P97 ; 3403P565
g3408P566 and 218P91 242P97 ; 3408P566
g3413P567 and 226P93 242P97 ; 3413P567
g3418P568 and 234P95 242P97 ; 3418P568
g2758P569 and 241P96 335P123 ; 2758P569
g2760P575 and 233P94 335P123 ; 2760P575
g2762P581 and 225P92 335P123 ; 2762P581
g2764P587 and 217P90 335P123 ; 2764P587
g2766P593 and 209P88 335P123 ; 2766P593
g1668P599 and 185P80 1689P157 1690P158 ; 1668P599
g2339P600 and 185P80 1691P159 1694P160 ; 2339P600
g1661P601 and 179P78 1689P157 1690P158 ; 1661P601
g2332P602 and 179P78 1691P159 1694P160 ; 2332P602
g2260P603 and 173P76 1691P159 1694P160 ; 2260P603
g1586P604 and 173P76 1689P157 1690P158 ; 1586P604
g1580P605 and 170P75 1689P157 1690P158 ; 1580P605
g2254P606 and 170P75 1691P159 1694P160 ; 2254P606
g1592P607 and 167P74 1689P157 1690P158 ; 1592P607
g2266P608 and 167P74 1691P159 1694P160 ; 2266P608
g2272P609 and 164P73 1691P159 1694P160 ; 2272P609
g1598P610 and 164P73 1689P157 1690P158 ; 1598P610
g1604P611 and 161P72 1689P157 1690P158 ; 1604P611
g2278P612 and 161P72 1691P159 1694P160 ; 2278P612
g2345P613 and 158P71 1691P159 1694P160 ; 2345P613
g1674P614 and 158P71 1689P157 1690P158 ; 1674P614
g1680P615 and 152P69 1689P157 1690P158 ; 1680P615
g2351P616 and 152P69 1691P159 1694P160 ; 2351P616
g2357P617 and 146P67 1691P159 1694P160 ; 2357P617
g1686P618 and 146P67 1689P157 1690P158 ; 1686P618
g3724P170_b not 3724P170 ; 3724P170_b
g3734P629 and 123P53 3717P169 3724P170_b ; 3734P629
g3643P634 and 97P37 4092P176 ; 3643P634
g3637P635 and 97P37 4092P176 ; 3637P635
g3646P636 and 94P36 4092P176 ; 3646P636
g3640P637 and 94P36 4092P176 ; 3640P637
g2358P162_b not 2358P162 ; 2358P162_b
g3202P638 and 88P34 2358P162_b ; 3202P638
g3199P639 and 88P34 2358P162_b ; 3199P639
g3196P640 and 86P32 2358P162_b ; 3196P640
g3193P641 and 83P31 2358P162_b ; 3193P641
g210P89_b not 210P89 ; 210P89_b
g3548P166_b not 3548P166 ; 3548P166_b
g2592P666 and 210P89_b 3548P166_b ; 2592P666
g218P91_b not 218P91 ; 218P91_b
g2597P667 and 218P91_b 3548P166_b ; 2597P667
g226P93_b not 226P93 ; 226P93_b
g2602P668 and 226P93_b 3548P166_b ; 2602P668
g234P95_b not 234P95 ; 234P95_b
g2607P669 and 234P95_b 3548P166_b ; 2607P669
g257P102_b not 257P102 ; 257P102_b
g2686P670 and 257P102_b 3548P166_b ; 2686P670
g265P104_b not 265P104 ; 265P104_b
g2691P671 and 265P104_b 3548P166_b ; 2691P671
g273P106_b not 273P106 ; 273P106_b
g2696P672 and 273P106_b 3548P166_b ; 2696P672
g281P108_b not 281P108 ; 281P108_b
g2701P673 and 281P108_b 3548P166_b ; 2701P673
g324P120_b not 324P120 ; 324P120_b
g2996P674 and 324P120_b 3548P166_b ; 2996P674
g341P125_b not 341P125 ; 341P125_b
g3003P675 and 341P125_b 3548P166_b ; 3003P675
g351P127_b not 351P127 ; 351P127_b
g3008P676 and 351P127_b 3548P166_b ; 3008P676
g2869P677 and 2358P162 2822P361_b ; 2869P677
g2881P678 and 2358P162 2822P361_b ; 2881P678
g2877P679 and 2358P162 2822P361_b ; 2877P679
g2873P680 and 2358P162 2822P361_b ; 2873P680
g2868P681 and 2358P162_b 2822P361_b ; 2868P681
g2872P682 and 2358P162_b 2822P361_b ; 2872P682
g2876P683 and 2358P162_b 2822P361_b ; 2876P683
g2880P684 and 2358P162_b 2822P361_b ; 2880P684
g3239P685 and 251P100 351P127_b 534P149 ; 3239P685
g3550P167_b not 3550P167 ; 3550P167_b
g2990P686 and 351P127_b 534P149 3550P167_b ; 2990P686
g2984P687 and 341P125_b 523P148 3550P167_b ; 2984P687
g3235P688 and 251P100 341P125_b 523P148 ; 3235P688
g2975P691 and 324P120_b 503P146 3550P167_b ; 2975P691
g3229P692 and 251P100 324P120_b 503P146 ; 3229P692
g316P118_b not 316P118 ; 316P118_b
g3288P693 and 251P100 316P118_b 490P145 ; 3288P693
g2914P694 and 251P100 316P118_b 490P145 ; 2914P694
g308P116_b not 308P116 ; 308P116_b
g2910P695 and 251P100 308P116_b 479P144 ; 2910P695
g3284P696 and 251P100 308P116_b 479P144 ; 3284P696
g3391P697 and 218P91_b 251P100 468P143 ; 3391P697
g2574P698 and 218P91_b 468P143 3550P167_b ; 2574P698
g3387P699 and 210P89_b 251P100 457P142 ; 3387P699
g2568P700 and 210P89_b 457P142 3550P167_b ; 2568P700
g3336P701 and 206P87 248P99 446P141 ; 3336P701
g3329P702 and 206P87 248P99 446P141 ; 3329P702
g3399P703 and 234P95_b 251P100 435P140 ; 3399P703
g2586P704 and 234P95_b 435P140 3550P167_b ; 2586P704
g3395P705 and 226P93_b 251P100 422P139 ; 3395P705
g2580P706 and 226P93_b 422P139 3550P167_b ; 2580P706
g2674P707 and 273P106_b 411P138 3550P167_b ; 2674P707
g3065P708 and 251P100 273P106_b 411P138 ; 3065P708
g3061P709 and 251P100 265P104_b 400P137 ; 3061P709
g2668P710 and 265P104_b 400P137 3550P167_b ; 2668P710
g2662P711 and 257P102_b 389P136 3550P167_b ; 2662P711
g3057P712 and 251P100 257P102_b 389P136 ; 3057P712
g3069P713 and 251P100 281P108_b 374P134 ; 3069P713
g2680P714 and 281P108_b 374P134 3550P167_b ; 2680P714
g332P122_b not 332P122 ; 332P122_b
g3118P715 and 332P122_b 369P131 ; 3118P715
g369P131_b not 369P131 ; 369P131_b
g3422P716 or 361P129 369P131_b ; 3422P716
g3120P717 and 332P122_b 361P129 ; 3120P717
g361P129_b not 361P129 ; 361P129_b
g3423P718 or 361P129_b 369P131 ; 3423P718
g3122P719 and 332P122_b 351P127 ; 3122P719
g3431P720 or 341P125 351P127_b ; 3431P720
g3124P721 and 332P122_b 341P125 ; 3124P721
g3432P722 or 341P125_b 351P127 ; 3432P722
g3147P723 or 332P122_b 3126P492 ; 3147P723
g3127P724 and 324P120 332P122_b ; 3127P724
g3129P727 and 316P118 332P122_b ; 3129P727
g5106P728 or 308P116 316P118_b ; 5106P728
g5107P729 or 308P116_b 316P118 ; 5107P729
g3131P730 and 308P116 332P122_b ; 3131P730
g302P114_b not 302P114 ; 302P114_b
g5116P731 or 293P112 302P114_b ; 5116P731
g3133P732 and 302P114 332P122_b ; 3133P732
g293P112_b not 293P112 ; 293P112_b
g5117P735 or 293P112_b 302P114 ; 5117P735
g3135P736 and 293P112 332P122_b ; 3135P736
g335P123_b not 335P123 ; 335P123_b
g2747P737 and 289P110 335P123_b ; 2747P737
g289P110_b not 289P110 ; 289P110_b
g3895P738 or 281P108 289P110_b ; 3895P738
g2749P739 and 281P108 335P123_b ; 2749P739
g3896P740 or 281P108_b 289P110 ; 3896P740
g2751P741 and 273P106 335P123_b ; 2751P741
g3904P742 or 265P104 273P106_b ; 3904P742
g2753P743 and 265P104 335P123_b ; 2753P743
g3905P744 or 265P104_b 273P106 ; 3905P744
g3913P745 or 234P95 257P102_b ; 3913P745
g2755P746 and 257P102 335P123_b ; 2755P746
g2920P747 and 254P101 293P112_b ; 2920P747
g2924P748 and 254P101 308P116_b ; 2924P748
g2929P749 and 254P101 316P118_b ; 2929P749
g3075P750 and 254P101 257P102_b ; 3075P750
g3080P751 and 254P101 265P104_b ; 3080P751
g3085P752 and 254P101 273P106_b ; 3085P752
g3090P753 and 254P101 281P108_b ; 3090P753
g3405P754 and 210P89_b 254P101 ; 3405P754
g3410P755 and 218P91_b 254P101 ; 3410P755
g3415P756 and 226P93_b 254P101 ; 3415P756
g3420P757 and 234P95_b 254P101 ; 3420P757
g3244P758 and 254P101 324P120_b ; 3244P758
g3254P759 and 254P101 351P127_b ; 3254P759
g3250P760 and 254P101 341P125_b ; 3250P760
g3293P761 and 254P101 293P112_b ; 3293P761
g3300P762 and 254P101 316P118_b ; 3300P762
g3296P763 and 254P101 308P116_b ; 3296P763
g2907P764 and 251P100 302P114_b ; 2907P764
g3334P765 and 251P100 361P129_b ; 3334P765
g3327P766 and 251P100 361P129_b ; 3327P766
g3281P767 and 251P100 302P114_b ; 3281P767
g3341P768 and 206P87 242P97 ; 3341P768
g3345P769 and 206P87 242P97 ; 3345P769
g2757P770 and 234P95 335P123_b ; 2757P770
g3914P771 or 234P95_b 257P102 ; 3914P771
g5364P772 or 218P91 226P93_b ; 5364P772
g2759P773 and 226P93 335P123_b ; 2759P773
g2761P774 and 218P91 335P123_b ; 2761P774
g5365P775 or 218P91_b 226P93 ; 5365P775
g206P87_b not 206P87 ; 206P87_b
g5375P776 or 206P87_b 210P89 ; 5375P776
g2763P777 and 210P89 335P123_b ; 2763P777
g2765P783 and 206P87 335P123_b ; 2765P783
g1691P159_b not 1691P159 ; 1691P159_b
g2259P784 and 203P86 1691P159_b 1694P160 ; 2259P784
g1689P157_b not 1689P157 ; 1689P157_b
g1585P785 and 203P86 1689P157_b 1690P158 ; 1585P785
g2253P786 and 200P85 1691P159_b 1694P160 ; 2253P786
g1579P787 and 200P85 1689P157_b 1690P158 ; 1579P787
g2265P788 and 197P84 1691P159_b 1694P160 ; 2265P788
g1591P789 and 197P84 1689P157_b 1690P158 ; 1591P789
g2271P790 and 194P83 1691P159_b 1694P160 ; 2271P790
g1597P791 and 194P83 1689P157_b 1690P158 ; 1597P791
g2277P792 and 191P82 1691P159_b 1694P160 ; 2277P792
g1603P793 and 191P82 1689P157_b 1690P158 ; 1603P793
g1673P794 and 188P81 1689P157_b 1690P158 ; 1673P794
g2344P795 and 188P81 1691P159_b 1694P160 ; 2344P795
g2338P796 and 182P79 1691P159_b 1694P160 ; 2338P796
g1667P797 and 182P79 1689P157_b 1690P158 ; 1667P797
g2331P798 and 176P77 1691P159_b 1694P160 ; 2331P798
g1660P799 and 176P77 1689P157_b 1690P158 ; 1660P799
g2350P800 and 155P70 1691P159_b 1694P160 ; 2350P800
g1679P801 and 155P70 1689P157_b 1690P158 ; 1679P801
g1685P802 and 149P68 1689P157_b 1690P158 ; 1685P802
g2356P803 and 149P68 1691P159_b 1694P160 ; 2356P803
g3838P804 and 131P59 4091P175_b 4092P176 ; 3838P804
g3847P805 and 130P58 4091P175_b 4092P176 ; 3847P805
g3841P806 and 129P57 4091P175_b 4092P176 ; 3841P806
g3789P807 and 128P56 4091P175_b 4092P176 ; 3789P807
g3786P808 and 127P55 4091P175_b 4092P176 ; 3786P808
g3783P809 and 126P54 4091P175_b 4092P176 ; 3783P809
g4081P810 and 123P53 4091P175_b 4092P176 ; 4081P810
g4011P811 and 122P52 4091P175_b 4092P176 ; 4011P811
g4078P812 and 121P51 4091P175_b 4092P176 ; 4078P812
g3844P814 and 119P49 4091P175_b 4092P176 ; 3844P814
g3780P816 and 117P47 4091P175_b 4092P176 ; 3780P816
g4075P817 and 116P46 4091P175_b 4092P176 ; 4075P817
g4023P818 and 115P45 4091P175_b 4092P176 ; 4023P818
g4020P819 and 114P44 4091P175_b 4092P176 ; 4020P819
g4014P820 and 113P43 4091P175_b 4092P176 ; 4014P820
g4072P821 and 112P42 4091P175_b 4092P176 ; 4072P821
g3195P828 and 87P33 2358P162 ; 3195P828
g3192P829 and 83P31 2358P162 ; 3192P829
g4017P836 and 53P19 4091P175_b 4092P176 ; 4017P836
g4069P837 and 52P18 4091P175_b 4092P176 ; 4069P837
g3201P842 and 34P12 2358P162 ; 3201P842
g3198P843 and 34P12 2358P162 ; 3198P843
g3255P854 or 534P149 3253P480 3254P759 ; 3255P854
g3240P855 or 3238P409 3239P685 ; 3240P855
g3009P856 or 534P149 3006P396 3008P676 ; 3009P856
g2991P857 or 2988P410 2990P686 ; 2991P857
g2985P858 or 2982P413 2984P687 ; 2985P858
g3004P859 or 523P148 3001P395 3003P675 ; 3004P859
g3236P860 or 3234P414 3235P688 ; 3236P860
g3251P861 or 523P148 3249P486 3250P760 ; 3251P861
g3232P418_b not 3232P418 ; 3232P418_b
g5307P862 and 3247P417 3232P418_b ; 5307P862
g2979P420_b not 2979P420 ; 2979P420_b
g3015P863 and 2999P419 2979P420_b ; 3015P863
g2036P864 and 514P147 3147P723 ; 2036P864
g1789P865 and 514P147 3147P723 ; 1789P865
g2976P866 or 2973P423 2975P691 ; 2976P866
g2997P867 or 503P146 2994P394 2996P674 ; 2997P867
g3230P868 or 3228P424 3229P692 ; 3230P868
g3245P869 or 503P146 3243P498 3244P758 ; 3245P869
g3301P870 or 490P145 3299P507 3300P762 ; 3301P870
g3289P871 or 3287P427 3288P693 ; 3289P871
g2930P872 or 490P145 2927P510 2929P749 ; 2930P872
g2915P873 or 2913P428 2914P694 ; 2915P873
g2911P874 or 2909P431 2910P695 ; 2911P874
g2925P875 or 479P144 2922P518 2924P748 ; 2925P875
g3285P876 or 3283P432 3284P696 ; 3285P876
g3297P877 or 479P144 3295P515 3296P763 ; 3297P877
g3411P878 or 468P143 3408P566 3410P755 ; 3411P878
g3392P879 or 3390P435 3391P697 ; 3392P879
g2598P880 or 468P143 2595P387 2597P667 ; 2598P880
g2575P881 or 2572P436 2574P698 ; 2575P881
g3388P882 or 3386P439 3387P699 ; 3388P882
g3406P883 or 457P142 3403P565 3405P754 ; 3406P883
g2569P884 or 2566P440 2568P700 ; 2569P884
g2593P885 or 457P142 2590P386 2592P666 ; 2593P885
g3337P886 and 206P87_b 251P100 446P141 ; 3337P886
g3330P887 and 206P87_b 251P100 446P141 ; 3330P887
g3421P888 or 435P140 3418P568 3420P757 ; 3421P888
g3400P889 or 3398P445 3399P703 ; 3400P889
g2608P890 or 435P140 2605P389 2607P669 ; 2608P890
g2587P891 or 2584P446 2586P704 ; 2587P891
g3396P892 or 3394P449 3395P705 ; 3396P892
g3416P893 or 422P139 3413P567 3415P756 ; 3416P893
g2581P894 or 2578P450 2580P706 ; 2581P894
g2603P895 or 422P139 2600P388 2602P668 ; 2603P895
g2675P896 or 2672P453 2674P707 ; 2675P896
g2697P897 or 411P138 2694P392 2696P672 ; 2697P897
g3066P898 or 3064P454 3065P708 ; 3066P898
g3086P899 or 411P138 3083P545 3085P752 ; 3086P899
g3081P900 or 400P137 3078P553 3080P751 ; 3081P900
g3062P901 or 3060P457 3061P709 ; 3062P901
g2692P902 or 400P137 2689P391 2691P671 ; 2692P902
g2669P903 or 2666P458 2668P710 ; 2669P903
g2663P904 or 2660P461 2662P711 ; 2663P904
g2687P905 or 389P136 2684P390 2686P670 ; 2687P905
g3058P906 or 3056P462 3057P712 ; 3058P906
g3076P907 or 389P136 3073P560 3075P750 ; 3076P907
g3091P908 or 374P134 3088P539 3090P753 ; 3091P908
g3070P909 or 3068P466 3069P713 ; 3070P909
g2702P910 or 374P134 2699P393 2701P673 ; 2702P910
g2681P911 or 2678P467 2680P714 ; 2681P911
g5126P912 or 3119P470 3118P715 ; 5126P912
g3422P716_b not 3422P716 ; 3422P716_b
g3423P718_b not 3423P718 ; 3423P718_b
g3424P913 or 3422P716_b 3423P718_b ; 3424P913
g3137P914 or 3121P472 3120P717 ; 3137P914
g3335P915 or 3333P473 3334P765 ; 3335P915
g3328P916 or 3326P475 3327P766 ; 3328P916
g3139P917 or 3123P478 3122P719 ; 3139P917
g3431P720_b not 3431P720 ; 3431P720_b
g3432P722_b not 3432P722 ; 3432P722_b
g3433P918 or 3431P720_b 3432P722_b ; 3433P918
g3143P919 or 3125P485 3124P721 ; 3143P919
g3151P923 or 3128P497 3127P724 ; 3151P923
g3155P924 or 3130P505 3129P727 ; 3155P924
g5106P728_b not 5106P728 ; 5106P728_b
g5107P729_b not 5107P729 ; 5107P729_b
g5209P925 or 5106P728_b 5107P729_b ; 5209P925
g3161P926 or 3132P513 3131P730 ; 3161P926
g3165P927 or 3134P521 3133P732 ; 3165P927
g3282P928 or 3280P522 3281P767 ; 3282P928
g5116P731_b not 5116P731 ; 5116P731_b
g5117P735_b not 5117P735 ; 5117P735_b
g5206P929 or 5116P731_b 5117P735_b ; 5206P929
g2908P930 or 2906P525 2907P764 ; 2908P930
g3167P931 or 3136P529 3135P736 ; 3167P931
g5322P932 or 3292P531 3293P761 ; 5322P932
g2933P933 or 2918P533 2920P747 ; 2933P933
g5178P934 or 2748P535 2747P737 ; 5178P934
g3895P738_b not 3895P738 ; 3895P738_b
g3896P740_b not 3896P740 ; 3896P740_b
g3897P935 or 3895P738_b 3896P740_b ; 3897P935
g2767P936 or 2750P537 2749P739 ; 2767P936
g2772P937 or 2752P544 2751P741 ; 2772P937
g3904P742_b not 3904P742 ; 3904P742_b
g3905P744_b not 3905P744 ; 3905P744_b
g3906P938 or 3904P742_b 3905P744_b ; 3906P938
g2776P939 or 2754P551 2753P743 ; 2776P939
g2780P940 or 2756P558 2755P746 ; 2780P940
g3913P745_b not 3913P745 ; 3913P745_b
g3914P771_b not 3914P771 ; 3914P771_b
g3915P941 or 3913P745_b 3914P771_b ; 3915P941
g3342P942 and 206P87_b 254P101 ; 3342P942
g3346P943 and 206P87_b 254P101 ; 3346P943
g2784P944 or 2758P569 2757P770 ; 2784P944
g2788P945 or 2760P575 2759P773 ; 2788P945
g5364P772_b not 5364P772 ; 5364P772_b
g5365P775_b not 5365P775 ; 5365P775_b
g5399P946 or 5364P772_b 5365P775_b ; 5399P946
g2794P947 or 2762P581 2761P774 ; 2794P947
g2798P948 or 2764P587 2763P777 ; 2798P948
g5374P949 or 206P87 210P89_b ; 5374P949
g2802P950 or 2766P593 2765P783 ; 2802P950
g3203P951 or 3202P638 3201P842 ; 3203P951
g3200P952 or 3199P639 3198P843 ; 3200P952
g3197P953 or 3196P640 3195P828 ; 3197P953
g3194P954 or 3193P641 3192P829 ; 3194P954
g2870P955 and 82P30 2358P162_b 2822P361 ; 2870P955
g2875P956 and 81P29 2358P162 2822P361 ; 2875P956
g2871P957 and 80P28 2358P162 2822P361 ; 2871P957
g2866P958 and 79P27 2358P162_b 2822P361 ; 2866P958
g2874P959 and 26P9 2358P162_b 2822P361 ; 2874P959
g2879P960 and 25P8 2358P162 2822P361 ; 2879P960
g2878P961 and 24P7 2358P162_b 2822P361 ; 2878P961
g2867P962 and 23P6 2358P162 2822P361 ; 2867P962
g3845P963 and 4091P175_b 4092P176_b 3015P863 ; 3845P963
g2081P970 and 534P149 3139P917 ; 2081P970
g1823P971 and 534P149 3139P917 ; 1823P971
g1806P974 and 523P148 3143P919 ; 1806P974
g2059P975 and 523P148 3143P919 ; 2059P975
g3147P723_b not 3147P723 ; 3147P723_b
g2019P978 or 514P147 3147P723_b ; 2019P978
g1777P979 or 514P147 3147P723_b ; 1777P979
g2018P982 and 503P146 3151P923 ; 2018P982
g1775P983 and 503P146 3151P923 ; 1775P983
g490P145_b not 490P145 ; 490P145_b
g3155P924_b not 3155P924 ; 3155P924_b
g4812P986 and 490P145_b 3155P924_b ; 4812P986
g2001P987 and 490P145 3155P924 ; 2001P987
g1749P988 and 490P145 3155P924 ; 1749P988
g4716P989 and 490P145_b 3155P924_b ; 4716P989
g1742P992 and 479P144 3161P926 ; 1742P992
g1995P993 and 479P144 3161P926 ; 1995P993
g1064P996 and 468P143 2794P947 ; 1064P996
g1318P997 and 468P143 2794P947 ; 1318P997
g1301P1000 and 457P142 2798P948 ; 1301P1000
g1046P1001 and 457P142 2798P948 ; 1046P1001
g3347P1002 or 446P141 3345P769 3346P943 ; 3347P1002
g3338P1003 or 3336P701 3337P886 ; 3338P1003
g3343P1004 or 446P141 3341P768 3342P942 ; 3343P1004
g3331P1005 or 3329P702 3330P887 ; 3331P1005
g1031P1006 and 446P141 2802P950 ; 1031P1006
g1286P1007 and 446P141 2802P950 ; 1286P1007
g1341P1010 and 435P140 2784P944 ; 1341P1010
g1097P1011 and 435P140 2784P944 ; 1097P1011
g1071P1014 and 422P139 2788P945 ; 1071P1014
g422P139_b not 422P139 ; 422P139_b
g2788P945_b not 2788P945 ; 2788P945_b
g4228P1015 and 422P139_b 2788P945_b ; 4228P1015
g4348P1016 and 422P139_b 2788P945_b ; 4348P1016
g1324P1017 and 422P139 2788P945 ; 1324P1017
g1145P1020 and 411P138 2772P937 ; 1145P1020
g1404P1021 and 411P138 2772P937 ; 1404P1021
g1382P1024 and 400P137 2776P939 ; 1382P1024
g1128P1025 and 400P137 2776P939 ; 1128P1025
g1111P1028 and 389P136 2780P940 ; 1111P1028
g1359P1029 and 389P136 2780P940 ; 1359P1029
g374P134_b not 374P134 ; 374P134_b
g2767P936_b not 2767P936 ; 2767P936_b
g4464P1032 and 374P134_b 2767P936_b ; 4464P1032
g1412P1033 and 374P134 2767P936 ; 1412P1033
g1160P1034 and 374P134 2767P936 ; 1160P1034
g3514P1057 and 324P120_b 3424P913 3433P918 ; 3514P1057
g5375P776_b not 5375P776 ; 5375P776_b
g5374P949_b not 5374P949 ; 5374P949_b
g5396P1110 or 5375P776_b 5374P949_b ; 5396P1110
g2908P930_b not 2908P930 ; 2908P930_b
g4076P1118 and 4091P175_b 4092P176_b 2908P930_b ; 4076P1118
g4079P1119 and 4091P175_b 4092P176_b 2933P933 ; 4079P1119
g3335P915_b not 3335P915 ; 3335P915_b
g3836P1120 and 4091P175_b 4092P176_b 3335P915_b ; 3836P1120
g3717P169_b not 3717P169 ; 3717P169_b
g3731P1121 and 3717P169_b 3724P170_b 2933P933 ; 3731P1121
g3240P855_b not 3240P855 ; 3240P855_b
g5299P1122 and 3255P854 3240P855_b ; 5299P1122
g2991P857_b not 2991P857 ; 2991P857_b
g3021P1123 and 3009P856 2991P857_b ; 3021P1123
g3139P917_b not 3139P917 ; 3139P917_b
g2065P1124 or 534P149 3139P917_b ; 2065P1124
g1811P1125 or 534P149 3139P917_b ; 1811P1125
g2985P858_b not 2985P858 ; 2985P858_b
g3018P1126 and 2985P858_b 3004P859 ; 3018P1126
g3236P860_b not 3236P860 ; 3236P860_b
g5296P1127 and 3236P860_b 3251P861 ; 5296P1127
g3143P919_b not 3143P919 ; 3143P919_b
g1793P1128 or 523P148 3143P919_b ; 1793P1128
g2040P1129 or 523P148 3143P919_b ; 2040P1129
g514P147_b not 514P147 ; 514P147_b
g2020P1130 or 514P147_b 3147P723 ; 2020P1130
g1776P1131 or 514P147_b 3147P723 ; 1776P1131
g2976P866_b not 2976P866 ; 2976P866_b
g3012P1132 and 2976P866_b 2997P867 ; 3012P1132
g3230P868_b not 3230P868 ; 3230P868_b
g5304P1133 and 3230P868_b 3245P869 ; 5304P1133
g3151P923_b not 3151P923 ; 3151P923_b
g2007P1134 or 503P146 3151P923_b ; 2007P1134
g1766P1135 or 503P146 3151P923_b ; 1766P1135
g3289P871_b not 3289P871 ; 3289P871_b
g5315P1136 and 3301P870 3289P871_b ; 5315P1136
g2915P873_b not 2915P873 ; 2915P873_b
g2942P1137 and 2930P872 2915P873_b ; 2942P1137
g2097P1138 or 490P145 3155P924_b ; 2097P1138
g1757P1141 or 490P145 3155P924_b ; 1757P1141
g2911P874_b not 2911P874 ; 2911P874_b
g2939P1144 and 2911P874_b 2925P875 ; 2939P1144
g3285P876_b not 3285P876 ; 3285P876_b
g5312P1145 and 3285P876_b 3297P877 ; 5312P1145
g3161P926_b not 3161P926 ; 3161P926_b
g1729P1146 or 479P144 3161P926_b ; 1729P1146
g1846P1147 and 3165P927_b 3167P931_b 1742P992 ; 1846P1147
g1849P1148 and 3165P927_b 1742P992 ; 1849P1148
g1852P1149 and 3165P927_b 1742P992 ; 1852P1149
g1982P1150 or 479P144 3161P926_b ; 1982P1150
g2122P1151 and 3165P927_b 1995P993 ; 2122P1151
g2116P1152 and 3165P927_b 3167P931_b 1995P993 ; 2116P1152
g2119P1153 and 3165P927_b 1995P993 ; 2119P1153
g3392P879_b not 3392P879 ; 3392P879_b
g5276P1154 and 3411P878 3392P879_b ; 5276P1154
g2575P881_b not 2575P881 ; 2575P881_b
g2615P1155 and 2598P880 2575P881_b ; 2615P1155
g2794P947_b not 2794P947 ; 2794P947_b
g1051P1156 or 468P143 2794P947_b ; 1051P1156
g1305P1157 or 468P143 2794P947_b ; 1305P1157
g3388P882_b not 3388P882 ; 3388P882_b
g5289P1158 and 3388P882_b 3406P883 ; 5289P1158
g2569P884_b not 2569P884 ; 2569P884_b
g2611P1159 and 2569P884_b 2593P885 ; 2611P1159
g2798P948_b not 2798P948 ; 2798P948_b
g1287P1160 or 457P142 2798P948_b ; 1287P1160
g1033P1161 or 457P142 2798P948_b ; 1033P1161
g2802P950_b not 2802P950 ; 2802P950_b
g1022P1164 or 446P141 2802P950_b ; 1022P1164
g1276P1165 or 446P141 2802P950_b ; 1276P1165
g3400P889_b not 3400P889 ; 3400P889_b
g5268P1166 and 3421P888 3400P889_b ; 5268P1166
g2587P891_b not 2587P891 ; 2587P891_b
g2623P1167 and 2608P890 2587P891_b ; 2623P1167
g2784P944_b not 2784P944 ; 2784P944_b
g1330P1168 or 435P140 2784P944_b ; 1330P1168
g1088P1169 or 435P140 2784P944_b ; 1088P1169
g3396P892_b not 3396P892 ; 3396P892_b
g5279P1170 and 3396P892_b 3416P893 ; 5279P1170
g2581P894_b not 2581P894 ; 2581P894_b
g2619P1171 and 2581P894_b 2603P895 ; 2619P1171
g1079P1172 or 422P139 2788P945_b ; 1079P1172
g1420P1175 or 422P139 2788P945_b ; 1420P1175
g2675P896_b not 2675P896 ; 2675P896_b
g2713P1178 and 2675P896_b 2697P897 ; 2713P1178
g3066P898_b not 3066P898 ; 3066P898_b
g5263P1179 and 3066P898_b 3086P899 ; 5263P1179
g2772P937_b not 2772P937 ; 2772P937_b
g1133P1180 or 411P138 2772P937_b ; 1133P1180
g1388P1181 or 411P138 2772P937_b ; 1388P1181
g3062P901_b not 3062P901 ; 3062P901_b
g5260P1182 and 3081P900 3062P901_b ; 5260P1182
g2669P903_b not 2669P903 ; 2669P903_b
g2709P1183 and 2692P902 2669P903_b ; 2709P1183
g2776P939_b not 2776P939 ; 2776P939_b
g1363P1184 or 400P137 2776P939_b ; 1363P1184
g1115P1185 or 400P137 2776P939_b ; 1115P1185
g2663P904_b not 2663P904 ; 2663P904_b
g2705P1186 and 2663P904_b 2687P905 ; 2705P1186
g3058P906_b not 3058P906 ; 3058P906_b
g5271P1187 and 3058P906_b 3076P907 ; 5271P1187
g2780P940_b not 2780P940 ; 2780P940_b
g1099P1188 or 389P136 2780P940_b ; 1099P1188
g1342P1189 or 389P136 2780P940_b ; 1342P1189
g3070P909_b not 3070P909 ; 3070P909_b
g3852P1190 and 3091P908 3070P909_b ; 3852P1190
g2681P911_b not 2681P911 ; 2681P911_b
g2717P1191 and 2702P910 2681P911_b ; 2717P1191
g1428P1192 or 374P134 2767P936_b ; 1428P1192
g1151P1195 or 374P134 2767P936_b ; 1151P1195
g3452P1196 or 5126P912 3137P914_b ; 3452P1196
g3462P1210 or 3147P723 3151P923_b ; 3462P1210
g3424P913_b not 3424P913 ; 3424P913_b
g3433P918_b not 3433P918 ; 3433P918_b
g3517P1214 and 324P120_b 3424P913_b 3433P918_b ; 3517P1214
g3516P1215 and 324P120 3424P913 3433P918_b ; 3516P1215
g3513P1216 and 324P120 3424P913_b 3433P918 ; 3513P1216
g5209P925_b not 5209P925 ; 5209P925_b
g5214P1220 or 5209P925_b 5206P929 ; 5214P1220
g1845P1226 and 3165P927 3167P931_b ; 1845P1226
g2115P1229 and 3165P927 3167P931_b ; 2115P1229
g5330P1231 or 3282P928 5322P932 ; 5330P1231
g5206P929_b not 5206P929 ; 5206P929_b
g5215P1233 or 5209P925 5206P929_b ; 5215P1233
g3484P1241 or 5178P934 2802P950_b ; 3484P1241
g3955P1242 and 3897P935 3906P938 3915P941 ; 3955P1242
g3897P935_b not 3897P935 ; 3897P935_b
g3906P938_b not 3906P938 ; 3906P938_b
g3958P1243 and 3897P935_b 3906P938_b 3915P941 ; 3958P1243
g5396P1110_b not 5396P1110 ; 5396P1110_b
g5405P1264 or 5399P946 5396P1110_b ; 5405P1264
g1875P1279 and 54P20 3137P914_b ; 1875P1279
g4067P1284 and 4091P175_b 4092P176_b 3012P1132 ; 4067P1284
g4070P1285 and 4091P175_b 4092P176_b 2942P1137 ; 4070P1285
g4073P1286 and 4091P175_b 4092P176_b 2939P1144 ; 4073P1286
g4009P1287 and 4091P175_b 4092P176_b 2623P1167 ; 4009P1287
g4012P1288 and 4091P175_b 4092P176_b 2619P1171 ; 4012P1288
g4015P1289 and 4091P175_b 4092P176_b 2615P1155 ; 4015P1289
g4018P1290 and 4091P175_b 4092P176_b 2611P1159 ; 4018P1290
g3839P1291 and 4091P175_b 4092P176_b 3021P1123 ; 3839P1291
g3842P1292 and 4091P175_b 4092P176_b 3018P1126 ; 3842P1292
g3778P1293 and 4091P175_b 4092P176_b 2717P1191 ; 3778P1293
g3781P1294 and 4091P175_b 4092P176_b 2713P1178 ; 3781P1294
g3784P1295 and 4091P175_b 4092P176_b 2709P1183 ; 3784P1295
g3787P1296 and 4091P175_b 4092P176_b 2705P1186 ; 3787P1296
g534P149_b not 534P149 ; 534P149_b
g2066P1299 or 534P149_b 3139P917 ; 2066P1299
g1810P1300 or 534P149_b 3139P917 ; 1810P1300
g523P148_b not 523P148 ; 523P148_b
g1792P1303 or 523P148_b 3143P919 ; 1792P1303
g2041P1304 or 523P148_b 3143P919 ; 2041P1304
g5304P1133_b not 5304P1133 ; 5304P1133_b
g3891P1305 or 5307P862 5304P1133_b ; 3891P1305
g2019P978_b not 2019P978 ; 2019P978_b
g2020P1130_b not 2020P1130 ; 2020P1130_b
g2021P1306 or 2019P978_b 2020P1130_b ; 2021P1306
g1777P979_b not 1777P979 ; 1777P979_b
g1776P1131_b not 1776P1131 ; 1776P1131_b
g1778P1307 or 1777P979_b 1776P1131_b ; 1778P1307
g503P146_b not 503P146 ; 503P146_b
g2008P1310 or 503P146_b 3151P923 ; 2008P1310
g1765P1311 or 503P146_b 3151P923 ; 1765P1311
g2098P1314 or 490P145_b 3155P924 ; 2098P1314
g1756P1316 or 490P145_b 3155P924 ; 1756P1316
g479P144_b not 479P144 ; 479P144_b
g1728P1320 or 479P144_b 3161P926 ; 1728P1320
g1983P1321 or 479P144_b 3161P926 ; 1983P1321
g468P143_b not 468P143 ; 468P143_b
g1050P1324 or 468P143_b 2794P947 ; 1050P1324
g1306P1325 or 468P143_b 2794P947 ; 1306P1325
g457P142_b not 457P142 ; 457P142_b
g1288P1328 or 457P142_b 2798P948 ; 1288P1328
g1032P1329 or 457P142_b 2798P948 ; 1032P1329
g3338P1003_b not 3338P1003 ; 3338P1003_b
g3353P1330 and 3347P1002 3338P1003_b ; 3353P1330
g3331P1005_b not 3331P1005 ; 3331P1005_b
g3350P1331 and 3343P1004 3331P1005_b ; 3350P1331
g446P141_b not 446P141 ; 446P141_b
g1021P1332 or 446P141_b 2802P950 ; 1021P1332
g1277P1333 or 446P141_b 2802P950 ; 1277P1333
g435P140_b not 435P140 ; 435P140_b
g1331P1336 or 435P140_b 2784P944 ; 1331P1336
g1087P1337 or 435P140_b 2784P944 ; 1087P1337
g1078P1340 or 422P139_b 2788P945 ; 1078P1340
g1421P1342 or 422P139_b 2788P945 ; 1421P1342
g411P138_b not 411P138 ; 411P138_b
g1132P1346 or 411P138_b 2772P937 ; 1132P1346
g1389P1347 or 411P138_b 2772P937 ; 1389P1347
g400P137_b not 400P137 ; 400P137_b
g1364P1350 or 400P137_b 2776P939 ; 1364P1350
g1114P1351 or 400P137_b 2776P939 ; 1114P1351
g389P136_b not 389P136 ; 389P136_b
g1098P1354 or 389P136_b 2780P940 ; 1098P1354
g1343P1355 or 389P136_b 2780P940 ; 1343P1355
g1429P1358 or 374P134_b 2767P936 ; 1429P1358
g1150P1360 or 374P134_b 2767P936 ; 1150P1360
g5126P912_b not 5126P912 ; 5126P912_b
g3453P1361 or 5126P912_b 3137P914 ; 3453P1361
g4756P1363 or 3137P914 1875P1279 ; 4756P1363
g3444P1368 or 3139P917_b 3143P919 ; 3444P1368
g3443P1369 or 3139P917 3143P919_b ; 3443P1369
g3461P1370 or 3147P723_b 3151P923 ; 3461P1370
g3517P1214_b not 3517P1214 ; 3517P1214_b
g3516P1215_b not 3516P1215 ; 3516P1215_b
g3518P1371 and 3517P1214_b 3516P1215_b ; 3518P1371
g3514P1057_b not 3514P1057 ; 3514P1057_b
g3513P1216_b not 3513P1216 ; 3513P1216_b
g3515P1372 and 3514P1057_b 3513P1216_b ; 3515P1372
g5150P1373 or 3155P924_b 3161P926 ; 5150P1373
g5214P1220_b not 5214P1220 ; 5214P1220_b
g5215P1233_b not 5215P1233 ; 5215P1233_b
g5239P1374 or 5214P1220_b 5215P1233_b ; 5239P1374
g5151P1375 or 3155P924 3161P926_b ; 5151P1375
g5160P1380 or 3165P927_b 3167P931 ; 5160P1380
g5161P1385 or 3165P927 3167P931_b ; 5161P1385
g3282P928_b not 3282P928 ; 3282P928_b
g5322P932_b not 5322P932 ; 5322P932_b
g5331P1387 or 3282P928_b 5322P932_b ; 5331P1387
g5178P934_b not 5178P934 ; 5178P934_b
g3485P1388 or 5178P934_b 2802P950 ; 3485P1388
g3915P941_b not 3915P941 ; 3915P941_b
g3957P1389 and 3897P935 3906P938_b 3915P941_b ; 3957P1389
g5194P1390 or 2767P936_b 2772P937 ; 5194P1390
g5195P1391 or 2767P936 2772P937_b ; 5195P1391
g3954P1392 and 3897P935_b 3906P938 3915P941_b ; 3954P1392
g5204P1393 or 2776P939_b 2780P940 ; 5204P1393
g5205P1394 or 2776P939 2780P940_b ; 5205P1394
g3466P1395 or 2784P944_b 2788P945 ; 3466P1395
g3467P1396 or 2784P944 2788P945_b ; 3467P1396
g5399P946_b not 5399P946 ; 5399P946_b
g5404P1397 or 5399P946_b 5396P1110 ; 5404P1397
g3475P1398 or 2794P947_b 2798P948 ; 3475P1398
g3476P1399 or 2794P947 2798P948_b ; 3476P1399
g1876P1400 or 54P20 3137P914 ; 1876P1400
g4021P1401 and 4091P175_b 4092P176_b 3353P1330 ; 4021P1401
g5299P1122_b not 5299P1122 ; 5299P1122_b
g3881P1402 or 5299P1122_b 5296P1127 ; 3881P1402
g2065P1124_b not 2065P1124 ; 2065P1124_b
g2066P1299_b not 2066P1299 ; 2066P1299_b
g2067P1403 or 2065P1124_b 2066P1299_b ; 2067P1403
g1811P1125_b not 1811P1125 ; 1811P1125_b
g1810P1300_b not 1810P1300 ; 1810P1300_b
g1812P1404 or 1811P1125_b 1810P1300_b ; 1812P1404
g5296P1127_b not 5296P1127 ; 5296P1127_b
g3882P1405 or 5299P1122 5296P1127_b ; 3882P1405
g1793P1128_b not 1793P1128 ; 1793P1128_b
g1792P1303_b not 1792P1303 ; 1792P1303_b
g1794P1406 or 1793P1128_b 1792P1303_b ; 1794P1406
g1866P1407 and 1806P974 1778P1307 ; 1866P1407
g2040P1129_b not 2040P1129 ; 2040P1129_b
g2041P1304_b not 2041P1304 ; 2041P1304_b
g2042P1408 or 2040P1129_b 2041P1304_b ; 2042P1408
g2146P1409 and 2059P975 2021P1306 ; 2146P1409
g2142P1410 and 2059P975 2021P1306 ; 2142P1410
g5307P862_b not 5307P862 ; 5307P862_b
g3890P1411 or 5307P862_b 5304P1133 ; 3890P1411
g2007P1134_b not 2007P1134 ; 2007P1134_b
g2008P1310_b not 2008P1310 ; 2008P1310_b
g2009P1416 or 2007P1134_b 2008P1310_b ; 2009P1416
g1766P1135_b not 1766P1135 ; 1766P1135_b
g1765P1311_b not 1765P1311 ; 1765P1311_b
g1767P1417 or 1766P1135_b 1765P1311_b ; 1767P1417
g5315P1136_b not 5315P1136 ; 5315P1136_b
g5320P1418 or 5315P1136_b 5312P1145 ; 5320P1418
g2097P1138_b not 2097P1138 ; 2097P1138_b
g2098P1314_b not 2098P1314 ; 2098P1314_b
g2099P1419 or 2097P1138_b 2098P1314_b ; 2099P1419
g1757P1141_b not 1757P1141 ; 1757P1141_b
g1756P1316_b not 1756P1316 ; 1756P1316_b
g1758P1420 or 1757P1141_b 1756P1316_b ; 1758P1420
g5312P1145_b not 5312P1145 ; 5312P1145_b
g5321P1421 or 5315P1136 5312P1145_b ; 5321P1421
g1729P1146_b not 1729P1146 ; 1729P1146_b
g1728P1320_b not 1728P1320 ; 1728P1320_b
g1730P1422 or 1729P1146_b 1728P1320_b ; 1730P1422
g1982P1150_b not 1982P1150 ; 1982P1150_b
g1983P1321_b not 1983P1321 ; 1983P1321_b
g1984P1423 or 1982P1150_b 1983P1321_b ; 1984P1423
g5276P1154_b not 5276P1154 ; 5276P1154_b
g5285P1424 or 5276P1154_b 5279P1170 ; 5285P1424
g1051P1156_b not 1051P1156 ; 1051P1156_b
g1050P1324_b not 1050P1324 ; 1050P1324_b
g1052P1426 or 1051P1156_b 1050P1324_b ; 1052P1426
g1305P1157_b not 1305P1157 ; 1305P1157_b
g1306P1325_b not 1306P1325 ; 1306P1325_b
g1307P1427 or 1305P1157_b 1306P1325_b ; 1307P1427
g1287P1160_b not 1287P1160 ; 1287P1160_b
g1288P1328_b not 1288P1328 ; 1288P1328_b
g1289P1428 or 1287P1160_b 1288P1328_b ; 1289P1428
g1033P1161_b not 1033P1161 ; 1033P1161_b
g1032P1329_b not 1032P1329 ; 1032P1329_b
g1034P1429 or 1033P1161_b 1032P1329_b ; 1034P1429
g1022P1164_b not 1022P1164 ; 1022P1164_b
g1021P1332_b not 1021P1332 ; 1021P1332_b
g1023P1432 or 1022P1164_b 1021P1332_b ; 1023P1432
g1276P1165_b not 1276P1165 ; 1276P1165_b
g1277P1333_b not 1277P1333 ; 1277P1333_b
g1278P1433 or 1276P1165_b 1277P1333_b ; 1278P1433
g5268P1166_b not 5268P1166 ; 5268P1166_b
g3870P1434 or 5268P1166_b 5271P1187 ; 3870P1434
g1330P1168_b not 1330P1168 ; 1330P1168_b
g1331P1336_b not 1331P1336 ; 1331P1336_b
g1332P1435 or 1330P1168_b 1331P1336_b ; 1332P1435
g1088P1169_b not 1088P1169 ; 1088P1169_b
g1087P1337_b not 1087P1337 ; 1087P1337_b
g1089P1436 or 1088P1169_b 1087P1337_b ; 1089P1436
g5279P1170_b not 5279P1170 ; 5279P1170_b
g5284P1437 or 5276P1154 5279P1170_b ; 5284P1437
g1079P1172_b not 1079P1172 ; 1079P1172_b
g1078P1340_b not 1078P1340 ; 1078P1340_b
g1080P1438 or 1079P1172_b 1078P1340_b ; 1080P1438
g1420P1175_b not 1420P1175 ; 1420P1175_b
g1421P1342_b not 1421P1342 ; 1421P1342_b
g1422P1439 or 1420P1175_b 1421P1342_b ; 1422P1439
g5263P1179_b not 5263P1179 ; 5263P1179_b
g3860P1441 or 5263P1179_b 5260P1182 ; 3860P1441
g1133P1180_b not 1133P1180 ; 1133P1180_b
g1132P1346_b not 1132P1346 ; 1132P1346_b
g1134P1442 or 1133P1180_b 1132P1346_b ; 1134P1442
g1388P1181_b not 1388P1181 ; 1388P1181_b
g1389P1347_b not 1389P1347 ; 1389P1347_b
g1390P1443 or 1388P1181_b 1389P1347_b ; 1390P1443
g5260P1182_b not 5260P1182 ; 5260P1182_b
g3861P1444 or 5263P1179 5260P1182_b ; 3861P1444
g1363P1184_b not 1363P1184 ; 1363P1184_b
g1364P1350_b not 1364P1350 ; 1364P1350_b
g1365P1445 or 1363P1184_b 1364P1350_b ; 1365P1445
g1115P1185_b not 1115P1185 ; 1115P1185_b
g1114P1351_b not 1114P1351 ; 1114P1351_b
g1116P1446 or 1115P1185_b 1114P1351_b ; 1116P1446
g5271P1187_b not 5271P1187 ; 5271P1187_b
g3869P1447 or 5268P1166 5271P1187_b ; 3869P1447
g1099P1188_b not 1099P1188 ; 1099P1188_b
g1098P1354_b not 1098P1354 ; 1098P1354_b
g1100P1448 or 1099P1188_b 1098P1354_b ; 1100P1448
g1342P1189_b not 1342P1189 ; 1342P1189_b
g1343P1355_b not 1343P1355 ; 1343P1355_b
g1344P1449 or 1342P1189_b 1343P1355_b ; 1344P1449
g1428P1192_b not 1428P1192 ; 1428P1192_b
g1429P1358_b not 1429P1358 ; 1429P1358_b
g1430P1451 or 1428P1192_b 1429P1358_b ; 1430P1451
g1151P1195_b not 1151P1195 ; 1151P1195_b
g1150P1360_b not 1150P1360 ; 1150P1360_b
g1152P1452 or 1151P1195_b 1150P1360_b ; 1152P1452
g3452P1196_b not 3452P1196 ; 3452P1196_b
g3453P1361_b not 3453P1361 ; 3453P1361_b
g3454P1453 or 3452P1196_b 3453P1361_b ; 3454P1453
g3444P1368_b not 3444P1368 ; 3444P1368_b
g3443P1369_b not 3443P1369 ; 3443P1369_b
g3445P1455 or 3444P1368_b 3443P1369_b ; 3445P1455
g3462P1210_b not 3462P1210 ; 3462P1210_b
g3461P1370_b not 3461P1370 ; 3461P1370_b
g3463P1456 or 3462P1210_b 3461P1370_b ; 3463P1456
g3518P1371_b not 3518P1371 ; 3518P1371_b
g3515P1372_b not 3515P1372 ; 3515P1372_b
g5236P1457 or 3518P1371_b 3515P1372_b ; 5236P1457
g5150P1373_b not 5150P1373 ; 5150P1373_b
g5151P1375_b not 5151P1375 ; 5151P1375_b
g5219P1458 or 5150P1373_b 5151P1375_b ; 5219P1458
g5160P1380_b not 5160P1380 ; 5160P1380_b
g5161P1385_b not 5161P1385 ; 5161P1385_b
g5216P1460 or 5160P1380_b 5161P1385_b ; 5216P1460
g5330P1231_b not 5330P1231 ; 5330P1231_b
g5331P1387_b not 5331P1387 ; 5331P1387_b
g5386P1461 or 5330P1231_b 5331P1387_b ; 5386P1461
g3484P1241_b not 3484P1241 ; 3484P1241_b
g3485P1388_b not 3485P1388 ; 3485P1388_b
g3486P1464 or 3484P1241_b 3485P1388_b ; 3486P1464
g3955P1242_b not 3955P1242 ; 3955P1242_b
g3954P1392_b not 3954P1392 ; 3954P1392_b
g3956P1465 and 3955P1242_b 3954P1392_b ; 3956P1465
g3958P1243_b not 3958P1243 ; 3958P1243_b
g3957P1389_b not 3957P1389 ; 3957P1389_b
g3959P1466 and 3958P1243_b 3957P1389_b ; 3959P1466
g5194P1390_b not 5194P1390 ; 5194P1390_b
g5195P1391_b not 5195P1391 ; 5195P1391_b
g5229P1467 or 5194P1390_b 5195P1391_b ; 5229P1467
g5204P1393_b not 5204P1393 ; 5204P1393_b
g5205P1394_b not 5205P1394 ; 5205P1394_b
g5226P1468 or 5204P1393_b 5205P1394_b ; 5226P1468
g3466P1395_b not 3466P1395 ; 3466P1395_b
g3467P1396_b not 3467P1396 ; 3467P1396_b
g3468P1469 or 3466P1395_b 3467P1396_b ; 3468P1469
g5405P1264_b not 5405P1264 ; 5405P1264_b
g5404P1397_b not 5404P1397 ; 5404P1397_b
g5425P1470 or 5405P1264_b 5404P1397_b ; 5425P1470
g3475P1398_b not 3475P1398 ; 3475P1398_b
g3476P1399_b not 3476P1399 ; 3476P1399_b
g3477P1471 or 3475P1398_b 3476P1399_b ; 3477P1471
g54P20_b not 54P20 ; 54P20_b
g1877P1472 or 54P20_b 3137P914_b ; 1877P1472
g3881P1402_b not 3881P1402 ; 3881P1402_b
g3882P1405_b not 3882P1405 ; 3882P1405_b
g3883P1473 or 3881P1402_b 3882P1405_b ; 3883P1473
g2147P1476 and 2081P970 2021P1306 2042P1408 ; 2147P1476
g2143P1477 and 2081P970 2021P1306 2042P1408 ; 2143P1477
g2133P1478 and 2081P970 2021P1306 2042P1408 2009P1416 ; 2133P1478
g2152P1479 and 2081P970 2042P1408 ; 2152P1479
g2149P1480 and 2081P970 2042P1408 ; 2149P1480
g1867P1481 and 1823P971 1778P1307 1794P1406 ; 1867P1481
g1861P1482 and 1823P971 1778P1307 1794P1406 1767P1417 ; 1861P1482
g1870P1483 and 1823P971 1794P1406 ; 1870P1483
g1860P1486 and 1806P974 1778P1307 1767P1417 ; 1860P1486
g2132P1489 and 2059P975 2021P1306 2009P1416 ; 2132P1489
g3891P1305_b not 3891P1305 ; 3891P1305_b
g3890P1411_b not 3890P1411 ; 3890P1411_b
g3892P1490 or 3891P1305_b 3890P1411_b ; 3892P1490
g2131P1493 and 2036P864 2009P1416 ; 2131P1493
g1859P1495 and 1789P865 1767P1417 ; 1859P1495
g5320P1418_b not 5320P1418 ; 5320P1418_b
g5321P1421_b not 5321P1421 ; 5321P1421_b
g5389P1499 or 5320P1418_b 5321P1421_b ; 5389P1499
g2158P1501 and 2099P1419 1984P1423 ; 2158P1501
g2120P1503 and 3165P927_b 2001P987 1984P1423 ; 2120P1503
g2117P1504 and 3165P927_b 3167P931_b 2001P987 1984P1423 ; 2117P1504
g2123P1505 and 3165P927_b 2001P987 1984P1423 ; 2123P1505
g2124P1506 and 2001P987 1984P1423 ; 2124P1506
g1855P1507 and 1758P1420 1730P1422 ; 1855P1507
g1847P1509 and 3165P927_b 3167P931_b 1749P988 1730P1422 ; 1847P1509
g1853P1510 and 3165P927_b 1749P988 1730P1422 ; 1853P1510
g1850P1511 and 3165P927_b 1749P988 1730P1422 ; 1850P1511
g1854P1512 and 1749P988 1730P1422 ; 1854P1512
g1856P1513 and 1749P988 1730P1422 ; 1856P1513
g5285P1424_b not 5285P1424 ; 5285P1424_b
g5284P1437_b not 5284P1437 ; 5284P1437_b
g5379P1518 or 5285P1424_b 5284P1437_b ; 5379P1518
g1173P1523 and 1052P1426 1034P1429 1080P1438 ; 1173P1523
g1177P1524 and 1052P1426 1080P1438 ; 1177P1524
g1169P1525 and 1064P996 1034P1429 1023P1432 ; 1169P1525
g1171P1526 and 1064P996 1034P1429 ; 1171P1526
g1174P1527 and 1064P996 1034P1429 ; 1174P1527
g1481P1528 and 1307P1427 1422P1439 ; 1481P1528
g1444P1531 and 1307P1427 1289P1428 1422P1439 ; 1444P1531
g1445P1533 and 1318P997 1289P1428 ; 1445P1533
g1440P1534 and 1318P997 1289P1428 1278P1433 ; 1440P1534
g1442P1535 and 1318P997 1289P1428 ; 1442P1535
g5295P1536 or 5289P1158 3350P1331_b ; 5295P1536
g1439P1539 and 1301P1000 1278P1433 ; 1439P1539
g1168P1542 and 1046P1001 1023P1432 ; 1168P1542
g3870P1434_b not 3870P1434 ; 3870P1434_b
g3869P1447_b not 3869P1447 ; 3869P1447_b
g3871P1548 or 3870P1434_b 3869P1447_b ; 3871P1548
g1170P1555 and 1071P1014 1052P1426 1034P1429 1023P1432 ; 1170P1555
g1175P1556 and 1071P1014 1052P1426 1034P1429 ; 1175P1556
g1172P1557 and 1071P1014 1052P1426 1034P1429 ; 1172P1557
g1176P1558 and 1071P1014 1052P1426 ; 1176P1558
g1178P1559 and 1071P1014 1052P1426 ; 1178P1559
g1443P1562 and 1324P1017 1307P1427 1289P1428 ; 1443P1562
g1441P1563 and 1324P1017 1307P1427 1289P1428 1278P1433 ; 1441P1563
g1446P1564 and 1324P1017 1307P1427 1289P1428 ; 1446P1564
g1447P1565 and 1324P1017 1307P1427 ; 1447P1565
g3860P1441_b not 3860P1441 ; 3860P1441_b
g3861P1444_b not 3861P1444 ; 3861P1444_b
g3862P1566 or 3860P1441_b 3861P1444_b ; 3862P1566
g1189P1567 and 1145P1020 1116P1446 1100P1448 ; 1189P1567
g1183P1568 and 1145P1020 1089P1436 1116P1446 1100P1448 ; 1183P1568
g1192P1569 and 1145P1020 1116P1446 ; 1192P1569
g1468P1572 and 1390P1443 1365P1445 1344P1449 1430P1451 ; 1468P1572
g1474P1573 and 1390P1443 1365P1445 1430P1451 ; 1474P1573
g1482P1575 and 1390P1443 1430P1451 ; 1482P1575
g1470P1576 and 1404P1021 1365P1445 1344P1449 ; 1470P1576
g1466P1577 and 1404P1021 1365P1445 1344P1449 ; 1466P1577
g1456P1578 and 1404P1021 1332P1435 1365P1445 1344P1449 ; 1456P1578
g1475P1579 and 1404P1021 1365P1445 ; 1475P1579
g1472P1580 and 1404P1021 1365P1445 ; 1472P1580
g1469P1583 and 1382P1024 1344P1449 ; 1469P1583
g1465P1584 and 1382P1024 1344P1449 ; 1465P1584
g1455P1585 and 1382P1024 1332P1435 1344P1449 ; 1455P1585
g1188P1587 and 1128P1025 1100P1448 ; 1188P1587
g1182P1588 and 1128P1025 1089P1436 1100P1448 ; 1182P1588
g1181P1590 and 1111P1028 1089P1436 ; 1181P1590
g1454P1593 and 1359P1029 1332P1435 ; 1454P1593
g1467P1596 and 1412P1033 1390P1443 1365P1445 1344P1449 ; 1467P1596
g1457P1597 and 1412P1033 1332P1435 1390P1443 1365P1445 1344P1449 ; 1457P1597
g1471P1598 and 1412P1033 1390P1443 1365P1445 1344P1449 ; 1471P1598
g1473P1599 and 1412P1033 1390P1443 1365P1445 ; 1473P1599
g1477P1600 and 1412P1033 1390P1443 ; 1477P1600
g1476P1601 and 1412P1033 1390P1443 1365P1445 ; 1476P1601
g1190P1603 and 1160P1034 1134P1442 1116P1446 1100P1448 ; 1190P1603
g1184P1604 and 1160P1034 1089P1436 1134P1442 1116P1446 1100P1448 ; 1184P1604
g1195P1605 and 1160P1034 1134P1442 ; 1195P1605
g1193P1606 and 1160P1034 1134P1442 1116P1446 ; 1193P1606
g1868P1609 and 3137P914 1778P1307 1812P1404 1794P1406 ; 1868P1609
g1862P1610 and 3137P914 1778P1307 1812P1404 1794P1406 1767P1417 ; 1862P1610
g1873P1611 and 3137P914 1812P1404 ; 1873P1611
g1871P1612 and 3137P914 1812P1404 1794P1406 ; 1871P1612
g2144P1613 and 3137P914 2021P1306 2067P1403 2042P1408 ; 2144P1613
g2134P1614 and 3137P914 2021P1306 2067P1403 2042P1408 2009P1416 ; 2134P1614
g2148P1615 and 3137P914 2021P1306 2067P1403 2042P1408 ; 2148P1615
g2150P1616 and 3137P914 2067P1403 2042P1408 ; 2150P1616
g2154P1617 and 3137P914 2067P1403 ; 2154P1617
g2153P1618 and 3137P914 2067P1403 2042P1408 ; 2153P1618
g2145P1620 and 3137P914_b 2021P1306 2067P1403 2042P1408 ; 2145P1620
g2159P1621 and 3137P914_b 2067P1403 ; 2159P1621
g2151P1622 and 3137P914_b 2067P1403 2042P1408 ; 2151P1622
g5236P1457_b not 5236P1457 ; 5236P1457_b
g3532P1627 or 5239P1374 5236P1457_b ; 3532P1627
g1851P1631 and 3165P927_b 1758P1420 1730P1422 ; 1851P1631
g2121P1633 and 3165P927_b 2099P1419 1984P1423 ; 2121P1633
g3956P1465_b not 3956P1465 ; 3956P1465_b
g3959P1466_b not 3959P1466 ; 3959P1466_b
g5422P1638 or 3956P1465_b 3959P1466_b ; 5422P1638
g132P60_b not 132P60 ; 132P60_b
g4107P1644 or 132P60_b 3167P931 ; 4107P1644
g1869P1645 and 54P20 3137P914_b 1778P1307 1812P1404 1794P1406 ; 1869P1645
g1874P1646 and 54P20 3137P914_b 1812P1404 ; 1874P1646
g1876P1400_b not 1876P1400 ; 1876P1400_b
g1877P1472_b not 1877P1472 ; 1877P1472_b
g1878P1647 or 1876P1400_b 1877P1472_b ; 1878P1647
g1872P1648 and 54P20 3137P914_b 1812P1404 1794P1406 ; 1872P1648
g1191P1649 and 4P1 1134P1442 1116P1446 1100P1448 1152P1452 ; 1191P1649
g1197P1650 and 4P1 1152P1452 ; 1197P1650
g1196P1651 and 4P1 1134P1442 1152P1452 ; 1196P1651
g1194P1652 and 4P1 1134P1442 1116P1446 1152P1452 ; 1194P1652
g3837P1653 and 4091P175 4092P176_b 1878P1647 ; 3837P1653
g2155P1657 or 2081P970 2154P1617 ; 2155P1657
g4748P1658 or 1823P971 1873P1611 1874P1646 ; 4748P1658
g4740P1661 or 1806P974 1870P1483 1871P1612 1872P1648 ; 4740P1661
g2059P975_b not 2059P975 ; 2059P975_b
g2152P1479_b not 2152P1479 ; 2152P1479_b
g2153P1618_b not 2153P1618 ; 2153P1618_b
g5009P1664 and 2059P975_b 2152P1479_b 2153P1618_b ; 5009P1664
g4928P1665 or 2059P975 2149P1480 2150P1616 2151P1622 ; 4928P1665
g2036P864_b not 2036P864 ; 2036P864_b
g2146P1409_b not 2146P1409 ; 2146P1409_b
g2147P1476_b not 2147P1476 ; 2147P1476_b
g2148P1615_b not 2148P1615 ; 2148P1615_b
g5029P1668 and 2036P864_b 2146P1409_b 2147P1476_b 2148P1615_b ; 5029P1668
g4941P1669 or 2036P864 2142P1410 2143P1477 2144P1613 2145P1620 ; 4941P1669
g4732P1670 or 1789P865 1866P1407 1867P1481 1868P1609 1869P1645 ; 4732P1670
g2135P1673 or 2018P982 2133P1478 2132P1489 2131P1493 2134P1614 ; 2135P1673
g1863P1675 or 1775P983 1861P1482 1860P1486 1859P1495 1862P1610 ; 1863P1675
g5389P1499_b not 5389P1499 ; 5389P1499_b
g5394P1676 or 5386P1461 5389P1499_b ; 5394P1676
g1730P1422_b not 1730P1422 ; 1730P1422_b
g1899P1680 or 1749P988 1730P1422_b ; 1899P1680
g1895P1681 or 4716P989 1730P1422_b ; 1895P1681
g1742P992_b not 1742P992 ; 1742P992_b
g1856P1513_b not 1856P1513 ; 1856P1513_b
g4708P1684 and 1742P992_b 1856P1513_b ; 4708P1684
g4700P1685 or 1742P992 1855P1507 1854P1512 ; 4700P1685
g2125P1688 or 1995P993 2124P1506 ; 2125P1688
g1064P996_b not 1064P996 ; 1064P996_b
g1178P1559_b not 1178P1559 ; 1178P1559_b
g4220P1693 and 1064P996_b 1178P1559_b ; 4220P1693
g4212P1694 or 1064P996 1177P1524 1176P1558 ; 4212P1694
g1448P1698 or 1318P997 1447P1565 ; 1448P1698
g5289P1158_b not 5289P1158 ; 5289P1158_b
g5294P1699 or 5289P1158_b 3350P1331 ; 5294P1699
g1301P1000_b not 1301P1000 ; 1301P1000_b
g1445P1533_b not 1445P1533 ; 1445P1533_b
g1446P1564_b not 1446P1564 ; 1446P1564_b
g4419P1702 and 1301P1000_b 1445P1533_b 1446P1564_b ; 4419P1702
g4361P1703 or 1301P1000 1444P1531 1442P1535 1443P1562 ; 4361P1703
g1046P1001_b not 1046P1001 ; 1046P1001_b
g1174P1527_b not 1174P1527 ; 1174P1527_b
g1175P1556_b not 1175P1556 ; 1175P1556_b
g4204P1706 and 1046P1001_b 1174P1527_b 1175P1556_b ; 4204P1706
g4196P1707 or 1046P1001 1173P1523 1171P1526 1172P1557 ; 4196P1707
g1458P1719 or 1341P1010 1456P1578 1455P1585 1454P1593 1457P1597 ; 1458P1719
g1185P1721 or 1097P1011 1183P1568 1182P1588 1181P1590 1184P1604 ; 1185P1721
g1052P1426_b not 1052P1426 ; 1052P1426_b
g1221P1722 or 1071P1014 1052P1426_b ; 1221P1722
g1217P1723 or 4228P1015 1052P1426_b ; 1217P1723
g4260P1727 or 1145P1020 1195P1605 1196P1651 ; 4260P1727
g1478P1731 or 1404P1021 1477P1600 ; 1478P1731
g1382P1024_b not 1382P1024 ; 1382P1024_b
g1475P1579_b not 1475P1579 ; 1475P1579_b
g1476P1601_b not 1476P1601 ; 1476P1601_b
g4555P1734 and 1382P1024_b 1475P1579_b 1476P1601_b ; 4555P1734
g4467P1735 or 1382P1024 1474P1573 1472P1580 1473P1599 ; 4467P1735
g4252P1737 or 1128P1025 1192P1569 1193P1606 1194P1652 ; 4252P1737
g4244P1739 or 1111P1028 1189P1567 1188P1587 1190P1603 1191P1649 ; 4244P1739
g1359P1029_b not 1359P1029 ; 1359P1029_b
g1470P1576_b not 1470P1576 ; 1470P1576_b
g1469P1583_b not 1469P1583 ; 1469P1583_b
g1471P1598_b not 1471P1598 ; 1471P1598_b
g4575P1742 and 1359P1029_b 1470P1576_b 1469P1583_b 1471P1598_b ; 4575P1742
g4487P1743 or 1359P1029 1468P1572 1466P1577 1465P1584 1467P1596 ; 4487P1743
g4268P1747 or 1160P1034 1197P1650 ; 4268P1747
g3520P1748 and 3454P1453 3445P1455 3463P1456 ; 3520P1748
g3454P1453_b not 3454P1453 ; 3454P1453_b
g3445P1455_b not 3445P1455 ; 3445P1455_b
g3523P1749 and 3454P1453_b 3445P1455_b 3463P1456 ; 3523P1749
g1812P1404_b not 1812P1404 ; 1812P1404_b
g1929P1751 or 4756P1363 1812P1404_b ; 1929P1751
g5219P1458_b not 5219P1458 ; 5219P1458_b
g5224P1756 or 5219P1458_b 5216P1460 ; 5224P1756
g5239P1374_b not 5239P1374 ; 5239P1374_b
g3531P1757 or 5239P1374_b 5236P1457 ; 3531P1757
g1852P1149_b not 1852P1149 ; 1852P1149_b
g1853P1510_b not 1853P1510 ; 1853P1510_b
g4692P1758 and 3165P927_b 1852P1149_b 1853P1510_b ; 4692P1758
g4684P1759 or 3165P927 1849P1148 1850P1511 1851P1631 ; 4684P1759
g2122P1151_b not 2122P1151 ; 2122P1151_b
g2123P1505_b not 2123P1505 ; 2123P1505_b
g4883P1760 and 3165P927_b 2122P1151_b 2123P1505_b ; 4883P1760
g4825P1761 or 3165P927 2119P1153 2120P1503 2121P1633 ; 4825P1761
g5216P1460_b not 5216P1460 ; 5216P1460_b
g5225P1762 or 5219P1458 5216P1460_b ; 5225P1762
g4111P1765 and 3167P931_b 4107P1644 ; 4111P1765
g3468P1469_b not 3468P1469 ; 3468P1469_b
g3477P1471_b not 3477P1471 ; 3477P1471_b
g3529P1767 and 3486P1464 3468P1469_b 3477P1471_b ; 3529P1767
g5422P1638_b not 5422P1638 ; 5422P1638_b
g3967P1769 or 5425P1470 5422P1638_b ; 3967P1769
g5229P1467_b not 5229P1467 ; 5229P1467_b
g5234P1771 or 5229P1467_b 5226P1468 ; 5234P1771
g5226P1468_b not 5226P1468 ; 5226P1468_b
g5235P1772 or 5229P1467 5226P1468_b ; 5235P1772
g3526P1773 and 3486P1464 3468P1469 3477P1471 ; 3526P1773
g4112P1774 and 132P60 4107P1644 ; 4112P1774
g1902P1775 and 54P20 1857P1608 ; 1902P1775
g1224P1777 and 4P1 1179P1552 ; 1224P1777
g1152P1452_b not 1152P1452 ; 1152P1452_b
g1198P1778 or 4P1 1152P1452_b ; 1198P1778
g4748P1658_b not 4748P1658 ; 4748P1658_b
g1925P1780 or 1794P1406 4748P1658_b ; 1925P1780
g4740P1661_b not 4740P1661 ; 4740P1661_b
g1920P1789 or 1778P1307 4740P1661_b ; 1920P1789
g4732P1670_b not 4732P1670 ; 4732P1670_b
g1915P1790 or 1767P1417 4732P1670_b ; 1915P1790
g1903P1793 or 1863P1675 1902P1775 ; 1903P1793
g4815P1794 or 2158P1501 2125P1688 ; 4815P1794
g1749P988_b not 1749P988 ; 1749P988_b
g1900P1795 or 1749P988_b 1730P1422 ; 1900P1795
g4716P989_b not 4716P989 ; 4716P989_b
g1896P1796 or 4716P989_b 1730P1422 ; 1896P1796
g4220P1693_b not 4220P1693 ; 4220P1693_b
g1214P1801 or 1034P1429 4220P1693_b ; 1214P1801
g4212P1694_b not 4212P1694 ; 4212P1694_b
g1211P1803 or 1034P1429 4212P1694_b ; 1211P1803
g4351P1805 or 1481P1528 1448P1698 ; 4351P1805
g5295P1536_b not 5295P1536 ; 5295P1536_b
g5294P1699_b not 5294P1699 ; 5294P1699_b
g5376P1808 or 5295P1536_b 5294P1699_b ; 5376P1808
g4204P1706_b not 4204P1706 ; 4204P1706_b
g1207P1811 or 1023P1432 4204P1706_b ; 1207P1811
g4196P1707_b not 4196P1707 ; 4196P1707_b
g1204P1813 or 1023P1432 4196P1707_b ; 1204P1813
g4244P1739_b not 4244P1739 ; 4244P1739_b
g1237P1818 or 1089P1436 4244P1739_b ; 1237P1818
g1225P1819 or 1185P1721 1224P1777 ; 1225P1819
g1071P1014_b not 1071P1014 ; 1071P1014_b
g1222P1820 or 1071P1014_b 1052P1426 ; 1222P1820
g4228P1015_b not 4228P1015 ; 4228P1015_b
g1218P1821 or 4228P1015_b 1052P1426 ; 1218P1821
g4260P1727_b not 4260P1727 ; 4260P1727_b
g1247P1822 or 1116P1446 4260P1727_b ; 1247P1822
g4268P1747_b not 4268P1747 ; 4268P1747_b
g1252P1824 or 1134P1442 4268P1747_b ; 1252P1824
g4477P1825 or 1482P1575 1478P1731 ; 4477P1825
g4252P1737_b not 4252P1737 ; 4252P1737_b
g1242P1829 or 1100P1448 4252P1737_b ; 1242P1829
g3852P1190_b not 3852P1190 ; 3852P1190_b
g3943P1834 and 3852P1190_b 3871P1548 3862P1566 ; 3943P1834
g3862P1566_b not 3862P1566 ; 3862P1566_b
g3946P1835 and 3852P1190 3871P1548 3862P1566_b ; 3946P1835
g4467P1735_b not 4467P1735 ; 4467P1735_b
g4472P1836 or 4464P1032 4467P1735_b ; 4472P1836
g4555P1734_b not 4555P1734 ; 4555P1734_b
g4560P1837 or 1412P1033 4555P1734_b ; 4560P1837
g3463P1456_b not 3463P1456 ; 3463P1456_b
g3519P1839 and 3454P1453 3445P1455_b 3463P1456_b ; 3519P1839
g4756P1363_b not 4756P1363 ; 4756P1363_b
g1930P1840 or 4756P1363_b 1812P1404 ; 1930P1840
g5009P1664_b not 5009P1664 ; 5009P1664_b
g5014P1841 or 3137P914 5009P1664_b ; 5014P1841
g4931P1842 or 2159P1621 2155P1657 ; 4931P1842
g3949P1843 and 3328P916 3883P1473 3892P1490 ; 3949P1843
g3328P916_b not 3328P916 ; 3328P916_b
g3883P1473_b not 3883P1473 ; 3883P1473_b
g3952P1844 and 3328P916_b 3883P1473_b 3892P1490 ; 3952P1844
g3522P1845 and 3454P1453_b 3445P1455 3463P1456_b ; 3522P1845
g5224P1756_b not 5224P1756 ; 5224P1756_b
g5225P1762_b not 5225P1762 ; 5225P1762_b
g5247P1847 or 5224P1756_b 5225P1762_b ; 5247P1847
g4708P1684_b not 4708P1684 ; 4708P1684_b
g1892P1848 or 3165P927_b 4708P1684_b ; 1892P1848
g4700P1685_b not 4700P1685 ; 4700P1685_b
g1889P1850 or 3165P927_b 4700P1685_b ; 1889P1850
g5386P1461_b not 5386P1461 ; 5386P1461_b
g5395P1856 or 5386P1461_b 5389P1499 ; 5395P1856
g4684P1759_b not 4684P1759 ; 4684P1759_b
g1882P1857 or 3167P931_b 4684P1759_b ; 1882P1857
g4692P1758_b not 4692P1758 ; 4692P1758_b
g1885P1858 or 3167P931_b 4692P1758_b ; 1885P1858
g4113P1859 or 4111P1765 4112P1774 ; 4113P1859
g5234P1771_b not 5234P1771 ; 5234P1771_b
g5235P1772_b not 5235P1772 ; 5235P1772_b
g5255P1860 or 5234P1771_b 5235P1772_b ; 5255P1860
g3486P1464_b not 3486P1464 ; 3486P1464_b
g3528P1861 and 3486P1464_b 3468P1469 3477P1471_b ; 3528P1861
g5425P1470_b not 5425P1470 ; 5425P1470_b
g3966P1862 or 5425P1470_b 5422P1638 ; 3966P1862
g3525P1863 and 3486P1464_b 3468P1469_b 3477P1471 ; 3525P1863
g4P1_b not 4P1 ; 4P1_b
g1199P1865 or 4P1_b 1152P1452 ; 1199P1865
g3733P1868 and 3717P169_b 3724P170 4113P1859 ; 3733P1868
g1694P160_b not 1694P160 ; 1694P160_b
g2335P1869 and 1691P159_b 1694P160_b 3848P1864 ; 2335P1869
g1690P158_b not 1690P158 ; 1690P158_b
g1664P1870 and 1689P157_b 1690P158_b 3848P1864 ; 1664P1870
g1794P1406_b not 1794P1406 ; 1794P1406_b
g1924P1872 or 1794P1406_b 4748P1658 ; 1924P1872
g4931P1842_b not 4931P1842 ; 4931P1842_b
g4936P1873 or 4928P1665 4931P1842_b ; 4936P1873
g1778P1307_b not 1778P1307 ; 1778P1307_b
g1919P1874 or 1778P1307_b 4740P1661 ; 1919P1874
g1767P1417_b not 1767P1417 ; 1767P1417_b
g1914P1875 or 1767P1417_b 4732P1670 ; 1914P1875
g5394P1676_b not 5394P1676 ; 5394P1676_b
g5395P1856_b not 5395P1856 ; 5395P1856_b
g5417P1877 or 5394P1676_b 5395P1856_b ; 5417P1877
g4815P1794_b not 4815P1794 ; 4815P1794_b
g4820P1879 or 4812P986 4815P1794_b ; 4820P1879
g4878P1880 or 2001P987 2125P1688 ; 4878P1880
g1758P1420_b not 1758P1420 ; 1758P1420_b
g1953P1881 and 1758P1420_b 1903P1793 ; 1953P1881
g1899P1680_b not 1899P1680 ; 1899P1680_b
g1900P1795_b not 1900P1795 ; 1900P1795_b
g1901P1882 or 1899P1680_b 1900P1795_b ; 1901P1882
g1895P1681_b not 1895P1681 ; 1895P1681_b
g1896P1796_b not 1896P1796 ; 1896P1796_b
g1897P1883 or 1895P1681_b 1896P1796_b ; 1897P1883
g5376P1808_b not 5376P1808 ; 5376P1808_b
g5385P1885 or 5379P1518 5376P1808_b ; 5385P1885
g1034P1429_b not 1034P1429 ; 1034P1429_b
g1213P1889 or 1034P1429_b 4220P1693 ; 1213P1889
g1210P1890 or 1034P1429_b 4212P1694 ; 1210P1890
g1023P1432_b not 1023P1432 ; 1023P1432_b
g1203P1891 or 1023P1432_b 4196P1707 ; 1203P1891
g1206P1892 or 1023P1432_b 4204P1706 ; 1206P1892
g1451P1551_b not 1451P1551 ; 1451P1551_b
g1458P1719_b not 1458P1719 ; 1458P1719_b
g1483P1895 and 1451P1551_b 1458P1719_b ; 1483P1895
g1089P1436_b not 1089P1436 ; 1089P1436_b
g1236P1896 or 1089P1436_b 4244P1739 ; 1236P1896
g1080P1438_b not 1080P1438 ; 1080P1438_b
g1272P1898 and 1080P1438_b 1225P1819 ; 1272P1898
g1221P1722_b not 1221P1722 ; 1221P1722_b
g1222P1820_b not 1222P1820 ; 1222P1820_b
g1223P1899 or 1221P1722_b 1222P1820_b ; 1223P1899
g1217P1723_b not 1217P1723 ; 1217P1723_b
g1218P1821_b not 1218P1821 ; 1218P1821_b
g1219P1900 or 1217P1723_b 1218P1821_b ; 1219P1900
g4351P1805_b not 4351P1805 ; 4351P1805_b
g4356P1901 or 4348P1016 4351P1805_b ; 4356P1901
g4414P1902 or 1324P1017 1448P1698 ; 4414P1902
g1134P1442_b not 1134P1442 ; 1134P1442_b
g1251P1903 or 1134P1442_b 4268P1747 ; 1251P1903
g1116P1446_b not 1116P1446 ; 1116P1446_b
g1246P1906 or 1116P1446_b 4260P1727 ; 1246P1906
g1100P1448_b not 1100P1448 ; 1100P1448_b
g1241P1907 or 1100P1448_b 4252P1737 ; 1241P1907
g3871P1548_b not 3871P1548 ; 3871P1548_b
g3945P1908 and 3852P1190_b 3871P1548_b 3862P1566_b ; 3945P1908
g3942P1909 and 3852P1190 3871P1548_b 3862P1566 ; 3942P1909
g4464P1032_b not 4464P1032 ; 4464P1032_b
g4473P1910 or 4464P1032_b 4467P1735 ; 4473P1910
g1412P1033_b not 1412P1033 ; 1412P1033_b
g4561P1911 or 1412P1033_b 4555P1734 ; 4561P1911
g3520P1748_b not 3520P1748 ; 3520P1748_b
g3519P1839_b not 3519P1839 ; 3519P1839_b
g3521P1912 and 3520P1748_b 3519P1839_b ; 3521P1912
g3523P1749_b not 3523P1749 ; 3523P1749_b
g3522P1845_b not 3522P1845 ; 3522P1845_b
g3524P1913 and 3523P1749_b 3522P1845_b ; 3524P1913
g1929P1751_b not 1929P1751 ; 1929P1751_b
g1930P1840_b not 1930P1840 ; 1930P1840_b
g1931P1914 or 1929P1751_b 1930P1840_b ; 1931P1914
g5015P1915 or 3137P914_b 5009P1664 ; 5015P1915
g2128P1619_b not 2128P1619 ; 2128P1619_b
g2135P1673_b not 2135P1673 ; 2135P1673_b
g2160P1916 and 2128P1619_b 2135P1673_b ; 2160P1916
g3892P1490_b not 3892P1490 ; 3892P1490_b
g3951P1918 and 3328P916 3883P1473_b 3892P1490_b ; 3951P1918
g3948P1919 and 3328P916_b 3883P1473 3892P1490_b ; 3948P1919
g1891P1923 or 3165P927 4708P1684 ; 1891P1923
g1888P1924 or 3165P927 4700P1685 ; 1888P1924
g1881P1927 or 3167P931 4684P1759 ; 1881P1927
g1884P1928 or 3167P931 4692P1758 ; 1884P1928
g3529P1767_b not 3529P1767 ; 3529P1767_b
g3528P1861_b not 3528P1861 ; 3528P1861_b
g3530P1929 and 3529P1767_b 3528P1861_b ; 3530P1929
g3526P1773_b not 3526P1773 ; 3526P1773_b
g3525P1863_b not 3525P1863 ; 3525P1863_b
g3527P1932 and 3526P1773_b 3525P1863_b ; 3527P1932
g1198P1778_b not 1198P1778 ; 1198P1778_b
g1199P1865_b not 1199P1865 ; 1199P1865_b
g1200P1934 or 1198P1778_b 1199P1865_b ; 1200P1934
g3840P1935 and 4091P175 4092P176_b 1931P1914 ; 3840P1935
g3779P1936 and 4091P175 4092P176_b 1200P1934 ; 3779P1936
g1925P1780_b not 1925P1780 ; 1925P1780_b
g1924P1872_b not 1924P1872 ; 1924P1872_b
g1926P1937 or 1925P1780_b 1924P1872_b ; 1926P1937
g4928P1665_b not 4928P1665 ; 4928P1665_b
g4937P1938 or 4928P1665_b 4931P1842 ; 4937P1938
g1920P1789_b not 1920P1789 ; 1920P1789_b
g1919P1874_b not 1919P1874 ; 1919P1874_b
g1921P1939 or 1920P1789_b 1919P1874_b ; 1921P1939
g1915P1790_b not 1915P1790 ; 1915P1790_b
g1914P1875_b not 1914P1875 ; 1914P1875_b
g1916P1940 or 1915P1790_b 1914P1875_b ; 1916P1940
g1903P1793_b not 1903P1793 ; 1903P1793_b
g1947P1941 and 1903P1793_b 1901P1882 ; 1947P1941
g4812P986_b not 4812P986 ; 4812P986_b
g4821P1943 or 4812P986_b 4815P1794 ; 4821P1943
g2001P987_b not 2001P987 ; 2001P987_b
g2125P1688_b not 2125P1688 ; 2125P1688_b
g4879P1944 or 2001P987_b 2125P1688_b ; 4879P1944
g1952P1945 and 1758P1420 1903P1793_b ; 1952P1945
g5379P1518_b not 5379P1518 ; 5379P1518_b
g5384P1947 or 5379P1518_b 5376P1808 ; 5384P1947
g1214P1801_b not 1214P1801 ; 1214P1801_b
g1213P1889_b not 1213P1889 ; 1213P1889_b
g1215P1948 or 1214P1801_b 1213P1889_b ; 1215P1948
g1211P1803_b not 1211P1803 ; 1211P1803_b
g1210P1890_b not 1210P1890 ; 1210P1890_b
g1212P1949 or 1211P1803_b 1210P1890_b ; 1212P1949
g1207P1811_b not 1207P1811 ; 1207P1811_b
g1206P1892_b not 1206P1892 ; 1206P1892_b
g1208P1950 or 1207P1811_b 1206P1892_b ; 1208P1950
g1204P1813_b not 1204P1813 ; 1204P1813_b
g1203P1891_b not 1203P1891 ; 1203P1891_b
g1205P1951 or 1204P1813_b 1203P1891_b ; 1205P1951
g1237P1818_b not 1237P1818 ; 1237P1818_b
g1236P1896_b not 1236P1896 ; 1236P1896_b
g1238P1953 or 1237P1818_b 1236P1896_b ; 1238P1953
g1225P1819_b not 1225P1819 ; 1225P1819_b
g1266P1954 and 1225P1819_b 1223P1899 ; 1266P1954
g1271P1955 and 1080P1438 1225P1819_b ; 1271P1955
g4348P1016_b not 4348P1016 ; 4348P1016_b
g4357P1957 or 4348P1016_b 4351P1805 ; 4357P1957
g1324P1017_b not 1324P1017 ; 1324P1017_b
g1448P1698_b not 1448P1698 ; 1448P1698_b
g4415P1958 or 1324P1017_b 1448P1698_b ; 4415P1958
g1247P1822_b not 1247P1822 ; 1247P1822_b
g1246P1906_b not 1246P1906 ; 1246P1906_b
g1248P1959 or 1247P1822_b 1246P1906_b ; 1248P1959
g1252P1824_b not 1252P1824 ; 1252P1824_b
g1251P1903_b not 1251P1903 ; 1251P1903_b
g1253P1960 or 1252P1824_b 1251P1903_b ; 1253P1960
g1242P1829_b not 1242P1829 ; 1242P1829_b
g1241P1907_b not 1241P1907 ; 1241P1907_b
g1243P1961 or 1242P1829_b 1241P1907_b ; 1243P1961
g3943P1834_b not 3943P1834 ; 3943P1834_b
g3942P1909_b not 3942P1909 ; 3942P1909_b
g3944P1962 and 3943P1834_b 3942P1909_b ; 3944P1962
g3946P1835_b not 3946P1835 ; 3946P1835_b
g3945P1908_b not 3945P1908 ; 3945P1908_b
g3947P1963 and 3946P1835_b 3945P1908_b ; 3947P1963
g4472P1836_b not 4472P1836 ; 4472P1836_b
g4473P1910_b not 4473P1910 ; 4473P1910_b
g4474P1964 or 4472P1836_b 4473P1910_b ; 4474P1964
g4560P1837_b not 4560P1837 ; 4560P1837_b
g4561P1911_b not 4561P1911 ; 4561P1911_b
g4562P1965 or 4560P1837_b 4561P1911_b ; 4562P1965
g3521P1912_b not 3521P1912 ; 3521P1912_b
g3524P1913_b not 3524P1913 ; 3524P1913_b
g5244P1966 or 3521P1912_b 3524P1913_b ; 5244P1966
g5014P1841_b not 5014P1841 ; 5014P1841_b
g5015P1915_b not 5015P1915 ; 5015P1915_b
g5016P1968 or 5014P1841_b 5015P1915_b ; 5016P1968
g3949P1843_b not 3949P1843 ; 3949P1843_b
g3948P1919_b not 3948P1919 ; 3948P1919_b
g3950P1970 and 3949P1843_b 3948P1919_b ; 3950P1970
g3952P1844_b not 3952P1844 ; 3952P1844_b
g3951P1918_b not 3951P1918 ; 3951P1918_b
g3953P1971 and 3952P1844_b 3951P1918_b ; 3953P1971
g1892P1848_b not 1892P1848 ; 1892P1848_b
g1891P1923_b not 1891P1923 ; 1891P1923_b
g1893P1972 or 1892P1848_b 1891P1923_b ; 1893P1972
g1889P1850_b not 1889P1850 ; 1889P1850_b
g1888P1924_b not 1888P1924 ; 1888P1924_b
g1890P1973 or 1889P1850_b 1888P1924_b ; 1890P1973
g1882P1857_b not 1882P1857 ; 1882P1857_b
g1881P1927_b not 1881P1927 ; 1881P1927_b
g1883P1974 or 1882P1857_b 1881P1927_b ; 1883P1974
g1885P1858_b not 1885P1858 ; 1885P1858_b
g1884P1928_b not 1884P1928 ; 1884P1928_b
g1886P1975 or 1885P1858_b 1884P1928_b ; 1886P1975
g3530P1929_b not 3530P1929 ; 3530P1929_b
g3527P1932_b not 3527P1932 ; 3527P1932_b
g5252P1976 or 3530P1929_b 3527P1932_b ; 5252P1976
g4068P1980 and 4091P175 4092P176_b 1916P1940 ; 4068P1980
g4010P1981 and 4091P175 4092P176_b 1238P1953 ; 4010P1981
g3846P1982 and 4091P175 4092P176_b 1921P1939 ; 3846P1982
g3843P1983 and 4091P175 4092P176_b 1926P1937 ; 3843P1983
g3788P1984 and 4091P175 4092P176_b 1243P1961 ; 3788P1984
g3785P1985 and 4091P175 4092P176_b 1248P1959 ; 3785P1985
g3782P1986 and 4091P175 4092P176_b 1253P1960 ; 3782P1986
g2155P1657_b not 2155P1657 ; 2155P1657_b
g5016P1968_b not 5016P1968 ; 5016P1968_b
g5025P1987 or 2155P1657_b 5016P1968_b ; 5025P1987
g4936P1873_b not 4936P1873 ; 4936P1873_b
g4937P1938_b not 4937P1938 ; 4937P1938_b
g4938P1989 or 4936P1873_b 4937P1938_b ; 4938P1989
g1943P1992 and 1903P1793 1890P1973 ; 1943P1992
g1897P1883_b not 1897P1883 ; 1897P1883_b
g1948P1993 and 1903P1793 1897P1883_b ; 1948P1993
g1935P1994 and 1903P1793 1883P1974 ; 1935P1994
g4820P1879_b not 4820P1879 ; 4820P1879_b
g4821P1943_b not 4821P1943 ; 4821P1943_b
g4822P1995 or 4820P1879_b 4821P1943_b ; 4822P1995
g4878P1880_b not 4878P1880 ; 4878P1880_b
g4879P1944_b not 4879P1944 ; 4879P1944_b
g4880P1996 or 4878P1880_b 4879P1944_b ; 4880P1996
g1954P1997 or 1953P1881 1952P1945 ; 1954P1997
g5385P1885_b not 5385P1885 ; 5385P1885_b
g5384P1947_b not 5384P1947 ; 5384P1947_b
g5409P1998 or 5385P1885_b 5384P1947_b ; 5409P1998
g1262P2002 and 1225P1819 1212P1949 ; 1262P2002
g1219P1900_b not 1219P1900 ; 1219P1900_b
g1267P2003 and 1225P1819 1219P1900_b ; 1267P2003
g1257P2004 and 1225P1819 1205P1951 ; 1257P2004
g1273P2005 or 1272P1898 1271P1955 ; 1273P2005
g4356P1901_b not 4356P1901 ; 4356P1901_b
g4357P1957_b not 4357P1957 ; 4357P1957_b
g4358P2006 or 4356P1901_b 4357P1957_b ; 4358P2006
g4414P1902_b not 4414P1902 ; 4414P1902_b
g4415P1958_b not 4415P1958 ; 4415P1958_b
g4416P2007 or 4414P1902_b 4415P1958_b ; 4416P2007
g4474P1964_b not 4474P1964 ; 4474P1964_b
g4483P2010 or 4477P1825 4474P1964_b ; 4483P2010
g1478P1731_b not 1478P1731 ; 1478P1731_b
g4562P1965_b not 4562P1965 ; 4562P1965_b
g4571P2011 or 1478P1731_b 4562P1965_b ; 4571P2011
g3944P1962_b not 3944P1962 ; 3944P1962_b
g3947P1963_b not 3947P1963 ; 3947P1963_b
g5406P2013 or 3944P1962_b 3947P1963_b ; 5406P2013
g3950P1970_b not 3950P1970 ; 3950P1970_b
g3953P1971_b not 3953P1971 ; 3953P1971_b
g5414P2018 or 3950P1970_b 3953P1971_b ; 5414P2018
g5244P1966_b not 5244P1966 ; 5244P1966_b
g3537P2019 or 5247P1847 5244P1966_b ; 3537P2019
g5252P1976_b not 5252P1976 ; 5252P1976_b
g3542P2023 or 5255P1860 5252P1976_b ; 3542P2023
g4071P2026 and 4091P175 4092P176_b 1954P1997 ; 4071P2026
g4013P2027 and 4091P175 4092P176_b 1273P2005 ; 4013P2027
g2341P2032 and 1691P159_b 1694P160_b 3849P2024 ; 2341P2032
g2337P2033 and 1691P159 1694P160_b 3790P2025 ; 2337P2033
g1670P2034 and 1689P157_b 1690P158_b 3849P2024 ; 1670P2034
g1666P2035 and 1689P157 1690P158_b 3790P2025 ; 1666P2035
g5024P2036 or 2155P1657 5016P1968 ; 5024P2036
g4938P1989_b not 4938P1989 ; 4938P1989_b
g4947P2038 or 4941P1669 4938P1989_b ; 4947P2038
g1886P1975_b not 1886P1975 ; 1886P1975_b
g1934P2039 and 1903P1793_b 1886P1975_b ; 1934P2039
g1949P2040 or 1947P1941 1948P1993 ; 1949P2040
g1893P1972_b not 1893P1972 ; 1893P1972_b
g1942P2041 and 1903P1793_b 1893P1972_b ; 1942P2041
g5414P2018_b not 5414P2018 ; 5414P2018_b
g3964P2042 or 5417P1877 5414P2018_b ; 3964P2042
g4416P2007_b not 4416P2007 ; 4416P2007_b
g4425P2047 or 4419P1702 4416P2007_b ; 4425P2047
g4358P2006_b not 4358P2006 ; 4358P2006_b
g4367P2048 or 4361P1703 4358P2006_b ; 4367P2048
g1208P1950_b not 1208P1950 ; 1208P1950_b
g1256P2049 and 1225P1819_b 1208P1950_b ; 1256P2049
g1268P2050 or 1266P1954 1267P2003 ; 1268P2050
g1215P1948_b not 1215P1948 ; 1215P1948_b
g1261P2051 and 1225P1819_b 1215P1948_b ; 1261P2051
g4477P1825_b not 4477P1825 ; 4477P1825_b
g4482P2055 or 4477P1825_b 4474P1964 ; 4482P2055
g4570P2056 or 1478P1731 4562P1965 ; 4570P2056
g5247P1847_b not 5247P1847 ; 5247P1847_b
g3536P2059 or 5247P1847_b 5244P1966 ; 3536P2059
g4880P1996_b not 4880P1996 ; 4880P1996_b
g4889P2060 or 4883P1760 4880P1996_b ; 4889P2060
g4822P1995_b not 4822P1995 ; 4822P1995_b
g4831P2061 or 4825P1761 4822P1995_b ; 4831P2061
g5255P1860_b not 5255P1860 ; 5255P1860_b
g3541P2062 or 5255P1860_b 5252P1976 ; 3541P2062
g4074P2072 and 4091P175 4092P176_b 1949P2040 ; 4074P2072
g4016P2073 and 4091P175 4092P176_b 1268P2050 ; 4016P2073
g2347P2088 and 1691P159_b 1694P160_b 3850P2069 ; 2347P2088
g2353P2089 and 1691P159_b 1694P160_b 3851P2063 ; 2353P2089
g2250P2090 and 1691P159_b 1694P160_b 4082P2071 ; 2250P2090
g2355P2091 and 1691P159 1694P160_b 3793P2065 ; 2355P2091
g2349P2092 and 1691P159 1694P160_b 3792P2066 ; 2349P2092
g2343P2093 and 1691P159 1694P160_b 3791P2067 ; 2343P2093
g2252P2094 and 1691P159 1694P160_b 4024P2068 ; 2252P2094
g1676P2095 and 1689P157_b 1690P158_b 3850P2069 ; 1676P2095
g1682P2096 and 1689P157_b 1690P158_b 3851P2063 ; 1682P2096
g1576P2097 and 1689P157_b 1690P158_b 4082P2071 ; 1576P2097
g1684P2098 and 1689P157 1690P158_b 3793P2065 ; 1684P2098
g1678P2099 and 1689P157 1690P158_b 3792P2066 ; 1678P2099
g1672P2100 and 1689P157 1690P158_b 3791P2067 ; 1672P2100
g1578P2101 and 1689P157 1690P158_b 4024P2068 ; 1578P2101
g5025P1987_b not 5025P1987 ; 5025P1987_b
g5024P2036_b not 5024P2036 ; 5024P2036_b
g5026P2102 or 5025P1987_b 5024P2036_b ; 5026P2102
g4941P1669_b not 4941P1669 ; 4941P1669_b
g4946P2103 or 4941P1669_b 4938P1989 ; 4946P2103
g1944P2104 or 1943P1992 1942P2041 ; 1944P2104
g5417P1877_b not 5417P1877 ; 5417P1877_b
g3963P2107 or 5417P1877_b 5414P2018 ; 3963P2107
g5409P1998_b not 5409P1998 ; 5409P1998_b
g3960P2108 or 5409P1998_b 5406P2013 ; 3960P2108
g4419P1702_b not 4419P1702 ; 4419P1702_b
g4424P2109 or 4419P1702_b 4416P2007 ; 4424P2109
g4361P1703_b not 4361P1703 ; 4361P1703_b
g4366P2110 or 4361P1703_b 4358P2006 ; 4366P2110
g1263P2111 or 1262P2002 1261P2051 ; 1263P2111
g1258P2112 or 1257P2004 1256P2049 ; 1258P2112
g4483P2010_b not 4483P2010 ; 4483P2010_b
g4482P2055_b not 4482P2055 ; 4482P2055_b
g4484P2114 or 4483P2010_b 4482P2055_b ; 4484P2114
g4571P2011_b not 4571P2011 ; 4571P2011_b
g4570P2056_b not 4570P2056 ; 4570P2056_b
g4572P2115 or 4571P2011_b 4570P2056_b ; 4572P2115
g5406P2013_b not 5406P2013 ; 5406P2013_b
g3961P2116 or 5409P1998 5406P2013_b ; 3961P2116
g4883P1760_b not 4883P1760 ; 4883P1760_b
g4888P2118 or 4883P1760_b 4880P1996 ; 4888P2118
g4825P1761_b not 4825P1761 ; 4825P1761_b
g4830P2119 or 4825P1761_b 4822P1995 ; 4830P2119
g4080P2134 and 4091P175 4092P176_b 1936P2105 ; 4080P2134
g4077P2135 and 4091P175 4092P176_b 1944P2104 ; 4077P2135
g4022P2136 and 4091P175 4092P176_b 1258P2112 ; 4022P2136
g4019P2137 and 4091P175 4092P176_b 1263P2111 ; 4019P2137
g3735P2142 and 3717P169 3724P170 1936P2105 ; 3735P2142
g2256P2143 and 1691P159_b 1694P160_b 4083P2130 ; 2256P2143
g2258P2144 and 1691P159 1694P160_b 4025P2129 ; 2258P2144
g1582P2145 and 1689P157_b 1690P158_b 4083P2130 ; 1582P2145
g1584P2146 and 1689P157 1690P158_b 4025P2129 ; 1584P2146
g5026P2102_b not 5026P2102 ; 5026P2102_b
g5035P2148 or 5029P1668 5026P2102_b ; 5035P2148
g4947P2038_b not 4947P2038 ; 4947P2038_b
g4946P2103_b not 4946P2103 ; 4946P2103_b
g4948P2149 or 4947P2038_b 4946P2103_b ; 4948P2149
g3964P2042_b not 3964P2042 ; 3964P2042_b
g3963P2107_b not 3963P2107 ; 3963P2107_b
g3965P2153 or 3964P2042_b 3963P2107_b ; 3965P2153
g3960P2108_b not 3960P2108 ; 3960P2108_b
g3961P2116_b not 3961P2116 ; 3961P2116_b
g3962P2154 or 3960P2108_b 3961P2116_b ; 3962P2154
g4425P2047_b not 4425P2047 ; 4425P2047_b
g4424P2109_b not 4424P2109 ; 4424P2109_b
g4426P2155 or 4425P2047_b 4424P2109_b ; 4426P2155
g4367P2048_b not 4367P2048 ; 4367P2048_b
g4366P2110_b not 4366P2110 ; 4366P2110_b
g4368P2156 or 4367P2048_b 4366P2110_b ; 4368P2156
g4572P2115_b not 4572P2115 ; 4572P2115_b
g4581P2161 or 4575P1742 4572P2115_b ; 4581P2161
g4484P2114_b not 4484P2114 ; 4484P2114_b
g4493P2162 or 4487P1743 4484P2114_b ; 4493P2162
g4889P2060_b not 4889P2060 ; 4889P2060_b
g4888P2118_b not 4888P2118 ; 4888P2118_b
g4890P2165 or 4889P2060_b 4888P2118_b ; 4890P2165
g4831P2061_b not 4831P2061 ; 4831P2061_b
g4830P2119_b not 4830P2119 ; 4830P2119_b
g4832P2166 or 4831P2061_b 4830P2119_b ; 4832P2166
g4113P1859_b not 4113P1859 ; 4113P1859_b
g4096P2167 or 1936P2105_b 4113P1859_b ; 4096P2167
g3648P2192 and 4091P175_b 3962P2154 ; 3648P2192
g3651P2193 and 4091P175_b 3965P2153 ; 3651P2193
g2262P2198 and 1691P159_b 1694P160_b 4084P2180 ; 2262P2198
g2264P2199 and 1691P159 1694P160_b 4026P2185 ; 2264P2199
g1588P2200 and 1689P157_b 1690P158_b 4084P2180 ; 1588P2200
g1590P2201 and 1689P157 1690P158_b 4026P2185 ; 1590P2201
g5029P1668_b not 5029P1668 ; 5029P1668_b
g5034P2203 or 5029P1668_b 5026P2102 ; 5034P2203
g4890P2165_b not 4890P2165 ; 4890P2165_b
g4899P2207 or 2099P1419 4890P2165_b ; 4899P2207
g4832P2166_b not 4832P2166 ; 4832P2166_b
g4841P2208 or 2099P1419 4832P2166_b ; 4841P2208
g4426P2155_b not 4426P2155 ; 4426P2155_b
g4435P2212 or 1422P1439 4426P2155_b ; 4435P2212
g4368P2156_b not 4368P2156 ; 4368P2156_b
g4377P2213 or 1422P1439 4368P2156_b ; 4377P2213
g4575P1742_b not 4575P1742 ; 4575P1742_b
g4580P2214 or 4575P1742_b 4572P2115 ; 4580P2214
g4487P1743_b not 4487P1743 ; 4487P1743_b
g4492P2215 or 4487P1743_b 4484P2114 ; 4492P2215
g4948P2149_b not 4948P2149 ; 4948P2149_b
g4957P2216 or 3137P914_b 4948P2149_b ; 4957P2216
g2268P2251 and 1691P159_b 1694P160_b 4085P2232 ; 2268P2251
g2274P2252 and 1691P159_b 1694P160_b 4086P2231 ; 2274P2252
g2276P2253 and 1691P159 1694P160_b 4028P2234 ; 2276P2253
g2270P2254 and 1691P159 1694P160_b 4027P2235 ; 2270P2254
g1594P2255 and 1689P157_b 1690P158_b 4085P2232 ; 1594P2255
g1600P2256 and 1689P157_b 1690P158_b 4086P2231 ; 1600P2256
g1602P2257 and 1689P157 1690P158_b 4028P2234 ; 1602P2257
g1596P2258 and 1689P157 1690P158_b 4027P2235 ; 1596P2258
g5035P2148_b not 5035P2148 ; 5035P2148_b
g5034P2203_b not 5034P2203 ; 5034P2203_b
g5036P2259 or 5035P2148_b 5034P2203_b ; 5036P2259
g2099P1419_b not 2099P1419 ; 2099P1419_b
g4898P2261 or 2099P1419_b 4890P2165 ; 4898P2261
g4840P2262 or 2099P1419_b 4832P2166 ; 4840P2262
g1422P1439_b not 1422P1439 ; 1422P1439_b
g4434P2263 or 1422P1439_b 4426P2155 ; 4434P2263
g4376P2264 or 1422P1439_b 4368P2156 ; 4376P2264
g4581P2161_b not 4581P2161 ; 4581P2161_b
g4580P2214_b not 4580P2214 ; 4580P2214_b
g4582P2265 or 4581P2161_b 4580P2214_b ; 4582P2265
g4493P2162_b not 4493P2162 ; 4493P2162_b
g4492P2215_b not 4492P2215 ; 4492P2215_b
g4494P2266 or 4493P2162_b 4492P2215_b ; 4494P2266
g4956P2267 or 3137P914 4948P2149 ; 4956P2267
g4899P2207_b not 4899P2207 ; 4899P2207_b
g4898P2261_b not 4898P2261 ; 4898P2261_b
g4900P2281 or 4899P2207_b 4898P2261_b ; 4900P2281
g4841P2208_b not 4841P2208 ; 4841P2208_b
g4840P2262_b not 4840P2262 ; 4840P2262_b
g4842P2282 or 4841P2208_b 4840P2262_b ; 4842P2282
g4435P2212_b not 4435P2212 ; 4435P2212_b
g4434P2263_b not 4434P2263 ; 4434P2263_b
g4436P2283 or 4435P2212_b 4434P2263_b ; 4436P2283
g4377P2213_b not 4377P2213 ; 4377P2213_b
g4376P2264_b not 4376P2264 ; 4376P2264_b
g4378P2284 or 4377P2213_b 4376P2264_b ; 4378P2284
g4582P2265_b not 4582P2265 ; 4582P2265_b
g4591P2287 or 1430P1451 4582P2265_b ; 4591P2287
g4494P2266_b not 4494P2266 ; 4494P2266_b
g4503P2288 or 1430P1451 4494P2266_b ; 4503P2288
g5036P2259_b not 5036P2259 ; 5036P2259_b
g5045P2289 or 3137P914_b 5036P2259_b ; 5045P2289
g4957P2216_b not 4957P2216 ; 4957P2216_b
g4956P2267_b not 4956P2267 ; 4956P2267_b
g4958P2290 or 4957P2216_b 4956P2267_b ; 4958P2290
g4958P2290_b not 4958P2290 ; 4958P2290_b
g4967P2301 or 2067P1403 4958P2290_b ; 4967P2301
g4842P2282_b not 4842P2282 ; 4842P2282_b
g4851P2304 or 1984P1423 4842P2282_b ; 4851P2304
g4900P2281_b not 4900P2281 ; 4900P2281_b
g4909P2305 or 1984P1423 4900P2281_b ; 4909P2305
g4378P2284_b not 4378P2284 ; 4378P2284_b
g4387P2306 or 1307P1427 4378P2284_b ; 4387P2306
g4436P2283_b not 4436P2283 ; 4436P2283_b
g4445P2307 or 1307P1427 4436P2283_b ; 4445P2307
g1430P1451_b not 1430P1451 ; 1430P1451_b
g4590P2310 or 1430P1451_b 4582P2265 ; 4590P2310
g4502P2311 or 1430P1451_b 4494P2266 ; 4502P2311
g5044P2312 or 3137P914 5036P2259 ; 5044P2312
g2067P1403_b not 2067P1403 ; 2067P1403_b
g4966P2318 or 2067P1403_b 4958P2290 ; 4966P2318
g1984P1423_b not 1984P1423 ; 1984P1423_b
g4850P2319 or 1984P1423_b 4842P2282 ; 4850P2319
g4908P2320 or 1984P1423_b 4900P2281 ; 4908P2320
g1307P1427_b not 1307P1427 ; 1307P1427_b
g4386P2321 or 1307P1427_b 4378P2284 ; 4386P2321
g4444P2322 or 1307P1427_b 4436P2283 ; 4444P2322
g4591P2287_b not 4591P2287 ; 4591P2287_b
g4590P2310_b not 4590P2310 ; 4590P2310_b
g4592P2323 or 4591P2287_b 4590P2310_b ; 4592P2323
g4503P2288_b not 4503P2288 ; 4503P2288_b
g4502P2311_b not 4502P2311 ; 4502P2311_b
g4504P2324 or 4503P2288_b 4502P2311_b ; 4504P2324
g5045P2289_b not 5045P2289 ; 5045P2289_b
g5044P2312_b not 5044P2312 ; 5044P2312_b
g5046P2325 or 5045P2289_b 5044P2312_b ; 5046P2325
g4967P2301_b not 4967P2301 ; 4967P2301_b
g4966P2318_b not 4966P2318 ; 4966P2318_b
g4968P2326 or 4967P2301_b 4966P2318_b ; 4968P2326
g5046P2325_b not 5046P2325 ; 5046P2325_b
g5055P2327 or 2067P1403 5046P2325_b ; 5055P2327
g4851P2304_b not 4851P2304 ; 4851P2304_b
g4850P2319_b not 4850P2319 ; 4850P2319_b
g4852P2328 or 4851P2304_b 4850P2319_b ; 4852P2328
g4909P2305_b not 4909P2305 ; 4909P2305_b
g4908P2320_b not 4908P2320 ; 4908P2320_b
g4910P2329 or 4909P2305_b 4908P2320_b ; 4910P2329
g4387P2306_b not 4387P2306 ; 4387P2306_b
g4386P2321_b not 4386P2321 ; 4386P2321_b
g4388P2330 or 4387P2306_b 4386P2321_b ; 4388P2330
g4445P2307_b not 4445P2307 ; 4445P2307_b
g4444P2322_b not 4444P2322 ; 4444P2322_b
g4446P2331 or 4445P2307_b 4444P2322_b ; 4446P2331
g4504P2324_b not 4504P2324 ; 4504P2324_b
g4513P2332 or 1390P1443 4504P2324_b ; 4513P2332
g4592P2323_b not 4592P2323 ; 4592P2323_b
g4601P2333 or 1390P1443 4592P2323_b ; 4601P2333
g5054P2338 or 2067P1403_b 5046P2325 ; 5054P2338
g4968P2326_b not 4968P2326 ; 4968P2326_b
g4977P2339 or 2009P1416 4968P2326_b ; 4977P2339
g4446P2331_b not 4446P2331 ; 4446P2331_b
g4455P2344 or 1278P1433 4446P2331_b ; 4455P2344
g4388P2330_b not 4388P2330 ; 4388P2330_b
g4397P2345 or 1278P1433 4388P2330_b ; 4397P2345
g1390P1443_b not 1390P1443 ; 1390P1443_b
g4512P2346 or 1390P1443_b 4504P2324 ; 4512P2346
g4600P2347 or 1390P1443_b 4592P2323 ; 4600P2347
g4910P2329_b not 4910P2329 ; 4910P2329_b
g4919P2348 or 3167P931_b 4910P2329_b ; 4919P2348
g4852P2328_b not 4852P2328 ; 4852P2328_b
g4861P2349 or 3167P931_b 4852P2328_b ; 4861P2349
g5055P2327_b not 5055P2327 ; 5055P2327_b
g5054P2338_b not 5054P2338 ; 5054P2338_b
g5056P2350 or 5055P2327_b 5054P2338_b ; 5056P2350
g2009P1416_b not 2009P1416 ; 2009P1416_b
g4976P2351 or 2009P1416_b 4968P2326 ; 4976P2351
g1278P1433_b not 1278P1433 ; 1278P1433_b
g4454P2352 or 1278P1433_b 4446P2331 ; 4454P2352
g4396P2353 or 1278P1433_b 4388P2330 ; 4396P2353
g4513P2332_b not 4513P2332 ; 4513P2332_b
g4512P2346_b not 4512P2346 ; 4512P2346_b
g4514P2354 or 4513P2332_b 4512P2346_b ; 4514P2354
g4601P2333_b not 4601P2333 ; 4601P2333_b
g4600P2347_b not 4600P2347 ; 4600P2347_b
g4602P2355 or 4601P2333_b 4600P2347_b ; 4602P2355
g4918P2356 or 3167P931 4910P2329 ; 4918P2356
g4860P2357 or 3167P931 4852P2328 ; 4860P2357
g5056P2350_b not 5056P2350 ; 5056P2350_b
g5065P2359 or 2009P1416 5056P2350_b ; 5065P2359
g4977P2339_b not 4977P2339 ; 4977P2339_b
g4976P2351_b not 4976P2351 ; 4976P2351_b
g4978P2360 or 4977P2339_b 4976P2351_b ; 4978P2360
g4455P2344_b not 4455P2344 ; 4455P2344_b
g4454P2352_b not 4454P2352 ; 4454P2352_b
g4456P2361 or 4455P2344_b 4454P2352_b ; 4456P2361
g4397P2345_b not 4397P2345 ; 4397P2345_b
g4396P2353_b not 4396P2353 ; 4396P2353_b
g4398P2362 or 4397P2345_b 4396P2353_b ; 4398P2362
g4602P2355_b not 4602P2355 ; 4602P2355_b
g4611P2363 or 1332P1435 4602P2355_b ; 4611P2363
g4514P2354_b not 4514P2354 ; 4514P2354_b
g4523P2364 or 1332P1435 4514P2354_b ; 4523P2364
g4919P2348_b not 4919P2348 ; 4919P2348_b
g4918P2356_b not 4918P2356 ; 4918P2356_b
g4920P2367 or 4919P2348_b 4918P2356_b ; 4920P2367
g4861P2349_b not 4861P2349 ; 4861P2349_b
g4860P2357_b not 4860P2357 ; 4860P2357_b
g4862P2368 or 4861P2349_b 4860P2357_b ; 4862P2368
g4978P2360_b not 4978P2360 ; 4978P2360_b
g4987P2369 or 2042P1408 4978P2360_b ; 4987P2369
g5064P2370 or 2009P1416_b 5056P2350 ; 5064P2370
g4398P2362_b not 4398P2362 ; 4398P2362_b
g1488P2372 or 1289P1428 4398P2362_b ; 1488P2372
g4456P2361_b not 4456P2361 ; 4456P2361_b
g1493P2373 or 1289P1428 4456P2361_b ; 1493P2373
g1332P1435_b not 1332P1435 ; 1332P1435_b
g4610P2376 or 1332P1435_b 4602P2355 ; 4610P2376
g4522P2377 or 1332P1435_b 4514P2354 ; 4522P2377
g4862P2368_b not 4862P2368 ; 4862P2368_b
g2165P2378 or 3165P927_b 4862P2368_b ; 2165P2378
g4920P2367_b not 4920P2367 ; 4920P2367_b
g2170P2379 or 3165P927_b 4920P2367_b ; 2170P2379
g2042P1408_b not 2042P1408 ; 2042P1408_b
g4986P2382 or 2042P1408_b 4978P2360 ; 4986P2382
g5065P2359_b not 5065P2359 ; 5065P2359_b
g5064P2370_b not 5064P2370 ; 5064P2370_b
g5066P2383 or 5065P2359_b 5064P2370_b ; 5066P2383
g1289P1428_b not 1289P1428 ; 1289P1428_b
g1487P2384 or 1289P1428_b 4398P2362 ; 1487P2384
g1492P2385 or 1289P1428_b 4456P2361 ; 1492P2385
g4611P2363_b not 4611P2363 ; 4611P2363_b
g4610P2376_b not 4610P2376 ; 4610P2376_b
g4612P2386 or 4611P2363_b 4610P2376_b ; 4612P2386
g4523P2364_b not 4523P2364 ; 4523P2364_b
g4522P2377_b not 4522P2377 ; 4522P2377_b
g4524P2387 or 4523P2364_b 4522P2377_b ; 4524P2387
g2164P2388 or 3165P927 4862P2368 ; 2164P2388
g2169P2389 or 3165P927 4920P2367 ; 2169P2389
g5066P2383_b not 5066P2383 ; 5066P2383_b
g4997P2390 or 2042P1408 5066P2383_b ; 4997P2390
g4987P2369_b not 4987P2369 ; 4987P2369_b
g4986P2382_b not 4986P2382 ; 4986P2382_b
g4988P2391 or 4987P2369_b 4986P2382_b ; 4988P2391
g1488P2372_b not 1488P2372 ; 1488P2372_b
g1487P2384_b not 1487P2384 ; 1487P2384_b
g1489P2393 or 1488P2372_b 1487P2384_b ; 1489P2393
g1493P2373_b not 1493P2373 ; 1493P2373_b
g1492P2385_b not 1492P2385 ; 1492P2385_b
g1494P2394 or 1493P2373_b 1492P2385_b ; 1494P2394
g4612P2386_b not 4612P2386 ; 4612P2386_b
g4543P2397 or 1365P1445 4612P2386_b ; 4543P2397
g4524P2387_b not 4524P2387 ; 4524P2387_b
g4533P2398 or 1365P1445 4524P2387_b ; 4533P2398
g2165P2378_b not 2165P2378 ; 2165P2378_b
g2164P2388_b not 2164P2388 ; 2164P2388_b
g2166P2399 or 2165P2378_b 2164P2388_b ; 2166P2399
g2170P2379_b not 2170P2379 ; 2170P2379_b
g2169P2389_b not 2169P2389 ; 2169P2389_b
g2171P2400 or 2170P2379_b 2169P2389_b ; 2171P2400
g2174P161_b not 2174P161 ; 2174P161_b
g2190P2401 and 2174P161_b 2135P1673_b 2171P2400 ; 2190P2401
g2191P2402 and 2174P161_b 2135P1673 2166P2399 ; 2191P2402
g2160P1916_b not 2160P1916 ; 2160P1916_b
g2193P2403 and 2174P161 2160P1916_b 2166P2399 ; 2193P2403
g2192P2404 and 2174P161 2160P1916 2171P2400 ; 2192P2404
g1497P156_b not 1497P156 ; 1497P156_b
g1513P2405 and 1497P156_b 1458P1719_b 1494P2394 ; 1513P2405
g1514P2406 and 1497P156_b 1458P1719 1489P2393 ; 1514P2406
g1483P1895_b not 1483P1895 ; 1483P1895_b
g1516P2407 and 1497P156 1483P1895_b 1489P2393 ; 1516P2407
g1515P2408 and 1497P156 1483P1895 1494P2394 ; 1515P2408
g4996P2409 or 2042P1408_b 5066P2383 ; 4996P2409
g4988P2391_b not 4988P2391 ; 4988P2391_b
g2184P2411 or 2021P1306 4988P2391_b ; 2184P2411
g1365P1445_b not 1365P1445 ; 1365P1445_b
g4542P2412 or 1365P1445_b 4612P2386 ; 4542P2412
g4532P2413 or 1365P1445_b 4524P2387 ; 4532P2413
g5074P2414 or 2190P2401 2191P2402 2193P2403 2192P2404 ; 5074P2414
g4620P2415 or 1513P2405 1514P2406 1516P2407 1515P2408 ; 4620P2415
g4997P2390_b not 4997P2390 ; 4997P2390_b
g4996P2409_b not 4996P2409 ; 4996P2409_b
g4998P2416 or 4997P2390_b 4996P2409_b ; 4998P2416
g2021P1306_b not 2021P1306 ; 2021P1306_b
g2183P2417 or 2021P1306_b 4988P2391 ; 2183P2417
g4543P2397_b not 4543P2397 ; 4543P2397_b
g4542P2412_b not 4542P2412 ; 4542P2412_b
g4544P2418 or 4543P2397_b 4542P2412_b ; 4544P2418
g4533P2398_b not 4533P2398 ; 4533P2398_b
g4532P2413_b not 4532P2413 ; 4532P2413_b
g4534P2419 or 4533P2398_b 4532P2413_b ; 4534P2419
g4998P2416_b not 4998P2416 ; 4998P2416_b
g2187P2423 or 2021P1306 4998P2416_b ; 2187P2423
g2184P2411_b not 2184P2411 ; 2184P2411_b
g2183P2417_b not 2183P2417 ; 2183P2417_b
g2185P2424 or 2184P2411_b 2183P2417_b ; 2185P2424
g4544P2418_b not 4544P2418 ; 4544P2418_b
g1510P2427 or 1344P1449 4544P2418_b ; 1510P2427
g4534P2419_b not 4534P2419 ; 4534P2419_b
g1507P2428 or 1344P1449 4534P2419_b ; 1507P2428
g2195P2429 and 2174P161 2185P2424 ; 2195P2429
g2186P2430 or 2021P1306_b 4998P2416 ; 2186P2430
g1344P1449_b not 1344P1449 ; 1344P1449_b
g1509P2431 or 1344P1449_b 4544P2418 ; 1509P2431
g1506P2432 or 1344P1449_b 4534P2419 ; 1506P2432
g2187P2423_b not 2187P2423 ; 2187P2423_b
g2186P2430_b not 2186P2430 ; 2186P2430_b
g2188P2433 or 2187P2423_b 2186P2430_b ; 2188P2433
g1510P2427_b not 1510P2427 ; 1510P2427_b
g1509P2431_b not 1509P2431 ; 1509P2431_b
g1511P2434 or 1510P2427_b 1509P2431_b ; 1511P2434
g1507P2428_b not 1507P2428 ; 1507P2428_b
g1506P2432_b not 1506P2432 ; 1506P2432_b
g1508P2435 or 1507P2428_b 1506P2432_b ; 1508P2435
g1518P2436 and 1497P156 1508P2435 ; 1518P2436
g2188P2433_b not 2188P2433 ; 2188P2433_b
g2194P2439 and 2174P161_b 2188P2433_b ; 2194P2439
g1511P2434_b not 1511P2434 ; 1511P2434_b
g1517P2440 and 1497P156_b 1511P2434_b ; 1517P2440
g5077P2441 or 2195P2429 2194P2439 ; 5077P2441
g4623P2442 or 1518P2436 1517P2440 ; 4623P2442
g5077P2441_b not 5077P2441 ; 5077P2441_b
g2196P2443 or 5074P2414 5077P2441_b ; 2196P2443
g4623P2442_b not 4623P2442 ; 4623P2442_b
g1519P2445 or 4620P2415 4623P2442_b ; 1519P2445
g5074P2414_b not 5074P2414 ; 5074P2414_b
g2197P2447 or 5074P2414_b 5077P2441 ; 2197P2447
g4620P2415_b not 4620P2415 ; 4620P2415_b
g1520P2448 or 4620P2415_b 4623P2442 ; 1520P2448
g2196P2443_b not 2196P2443 ; 2196P2443_b
g2197P2447_b not 2197P2447 ; 2197P2447_b
g2198P2449 or 2196P2443_b 2197P2447_b ; 2198P2449
g1519P2445_b not 1519P2445 ; 1519P2445_b
g1520P2448_b not 1520P2448 ; 1520P2448_b
g1521P2450 or 1519P2445_b 1520P2448_b ; 1521P2450
g2198P2449_b not 2198P2449 ; 2198P2449_b
g3652P2457 and 4091P175 2198P2449_b ; 3652P2457
g1521P2450_b not 1521P2450 ; 1521P2450_b
g3649P2458 and 4091P175 1521P2450_b ; 3649P2458
g3657P2459 or 3648P2192 3649P2458 ; 3657P2459
g3658P2460 or 3651P2193 3652P2457 ; 3658P2460
g3636P2461 and 4092P176_b 3657P2459 ; 3636P2461
g3642P2462 and 4092P176_b 3657P2459 ; 3642P2462
g3639P2463 and 4092P176_b 3658P2460 ; 3639P2463
g3645P2464 and 4092P176_b 3658P2460 ; 3645P2464
g3655P2465 or 3643P634 3642P2462 ; 3655P2465
g3653P2466 or 3637P635 3636P2461 ; 3653P2466
g3656P2467 or 3646P636 3645P2464 ; 3656P2467
g3654P2468 or 3640P637 3639P2463 ; 3654P2468
g2328P2473 and 1691P159_b 1694P160_b 3654P2468 ; 2328P2473
g2330P2474 and 1691P159 1694P160_b 3653P2466 ; 2330P2474
g1657P2475 and 1689P157_b 1690P158_b 3654P2468 ; 1657P2475
g1659P2476 and 1689P157 1690P158_b 3653P2466 ; 1659P2476
g1662P2477 or 1661P601 1660P799 1657P2475 1659P2476 ; 1662P2477
g2333P2478 or 2332P602 2331P798 2328P2473 2330P2474 ; 2333P2478
