name C3540.iscas
i 1(0)
i 13(1)
i 20(2)
i 33(3)
i 41(4)
i 45(5)
i 50(6)
i 58(7)
i 68(8)
i 77(9)
i 87(10)
i 97(11)
i 107(12)
i 116(13)
i 124(14)
i 125(15)
i 128(16)
i 132(17)
i 137(18)
i 143(19)
i 150(20)
i 159(21)
i 169(22)
i 179(23)
i 190(24)
i 200(25)
i 213(26)
i 222(27)
i 223(28)
i 226(29)
i 232(30)
i 238(31)
i 244(32)
i 250(33)
i 257(34)
i 264(35)
i 270(36)
i 274(37)
i 283(38)
i 294(39)
i 303(40)
i 311(41)
i 317(42)
i 322(43)
i 326(44)
i 329(45)
i 330(46)
i 343(47)
i 1698(48)
i 2897(49)

o 353(405)
o 355(399)
o 361(940)
o 358(1161)
o 351(1247)
o 372(1243)
o 369(1321)
o 399(1428)
o 364(1484)
o 396(1504)
o 384(1553)
o 367(1585)
o 387(1616)
o 393(1605)
o 390(1603)
o 378(1597)
o 375(1624)
o 381(1626)
o 407(1657)
o 409(1670)
o 405(1717)
o 402(1718)

g1 and 343(47) ; 2868(50)
g2 and 330(46) ; 3419(51)
g3 and 270(36) ; 2960(52)
g4 and 264(35) ; 2957(53)
g5 and 264(35)* 257(34)* ; 587(54)
g6 and 257(34) ; 2950(55)
g7 and 250(33) ; 2947(56)
g8 and 244(32) ; 2942(57)
g9 and 238(31) ; 2939(58)
g10 and 232(30) ; 2934(59)
g11 and 226(29) ; 2931(60)
g12 and 213(26) ; 2865(61)
g13 and 200(25) ; 1048(62)
g14 and 190(24) ; 1035(63)
g15 and 179(23) ; 2478(64)
g16 and 116(13) ; 540(65)
g17 and 116(13) ; 530(66)
g18 and 107(12) ; 907(67)
g19 and 107(12) ; 851(68)
g20 and 107(12) ; 526(69)
g21 and 107(12) ; 517(70)
g22 and 97(11) ; 3103(71)
g23 and 97(11) ; 3095(72)
g24 and 97(11) ; 848(73)
g25 and 97(11) ; 845(74)
g26 and 97(11) ; 513(75)
g27 and 97(11) ; 504(76)
g28 and 87(10) ; 842(77)
g29 and 87(10) ; 839(78)
g30 and 87(10) ; 501(79)
g31 and 87(10) ; 492(80)
g32 and 77(9) ; 483(81)
g33 and 77(9) ; 479(82)
g34 and 77(9) ; 476(83)
g35 and 68(8) ; 898(84)
g36 and 68(8) ; 836(85)
g37 and 68(8) ; 833(86)
g38 and 68(8) ; 467(87)
g39 and 68(8) ; 463(88)
g40 and 68(8) ; 460(89)
g41 and 58(7) ; 3087(90)
g42 and 58(7) ; 3079(91)
g43 and 58(7) ; 831(92)
g44 and 58(7) ; 828(93)
g45 and 58(7) ; 456(94)
g46 and 58(7) ; 447(95)
g47 and 50(6) ; 826(96)
g48 and 50(6) ; 3007(97)
g49 and 50(6) ; 442(98)
g50 and 50(6) ; 432(99)
g51 and 45(5) ; 802(100)
g52 and 45(5) ; 799(101)
g53 and 45(5)* 41(4)* ; 798(102)
g54 and 41(4) ; 791(103)
g55 and 33(3) ; 2051(104)
g56 and 33(3)* 1698(48)* ; 1699(105)
g57 and 33(3) ; 780(106)
g58 and 33(3) ; 776(107)
g59 and 33(3) ; 758(108)
g60 and 41(4) 33(3) ; 788(109)
g61 and 20(2) ; 1828(110)
g62 and 20(2) ; 1540(111)
g63 and 179(23) 20(2) ; 1051(112)
g64 and 200(25) 20(2) ; 1050(113)
g65 and 200(25) 20(2) ; 1049(114)
g66 and 20(2) ; 1032(115)
g67 and 20(2) ; 741(116)
g68 and 20(2) ; 732(117)
g69 and 20(2) ; 736(118)
g70 and 13(1) ; 724(119)
g71 and 13(1) ; 717(120)
g72 and 20(2) 13(1) ; 731(121)
g73 and 33(3) 20(2) 1(0) ; 1827(122)
g74 and 13(1) 1(0) ; 1826(123)
g75 and 1(0) ; 714(124)
g76 and 1(0) ; 890(125)
g77 and 1(0) ; 704(126)
g78 and 1(0) ; 707(127)
g79 and 2868(50)* 2865(61)* ; 2871(128)
g80 and 2868(50)* 2865(61)* ; 2874(129)
g81 and 3419(51) ; 3425(130)
g82 and 2960(52) ; 2964(131)
g83 and 530(66) 270(36) ; 552(132)
g84 and 2957(53) ; 2963(133)
g85 and 517(70) 264(35) ; 551(134)
g86 and 2950(55) ; 2954(135)
g87 and 504(76) 257(34) ; 550(136)
g88 and 587(54) 250(33) ; 588(137)
g89 and 2947(56) ; 2953(138)
g90 and 492(80) 250(33) ; 549(139)
g91 and 2942(57) ; 2946(140)
g92 and 483(81) 244(32) ; 548(141)
g93 and 2939(58) ; 2945(142)
g94 and 467(87) 238(31) ; 547(143)
g95 and 2934(59) ; 2938(144)
g96 and 447(95) 232(30) ; 546(145)
g97 and 2931(60) ; 2937(146)
g98 and 432(99) 226(29) ; 545(147)
g99 and 1035(63)* 1032(115)* ; 1038(148)
g100 and 1035(63)* 1032(115)* ; 1043(149)
g101 and 2478(64) ; 2481(150)
g102 and 169(22)* 1540(111)* ; 1541(151)
g103 and 540(65) ; 3040(152)
g104 and 907(67) ; 3098(153)
g105 and 907(67) ; 3106(154)
g106 and 851(68) 848(73) 842(77) ; 905(155)
g107 and 851(68) 848(73) 842(77) ; 906(156)
g108 and 526(69) ; 3037(157)
g109 and 526(69) 513(75) ; 626(158)
g110 and 3103(71) ; 3109(159)
g111 and 3095(72) ; 3101(160)
g112 and 513(75) ; 3030(161)
g113 and 501(79) ; 3027(162)
g114 and 479(82) ; 3020(163)
g115 and 476(83) 460(89) ; 635(164)
g116 and 898(84) ; 3082(165)
g117 and 898(84) ; 3090(166)
g118 and 836(85) 831(92) 826(96) ; 625(167)
g119 and 836(85) 831(92) 826(96) ; 897(168)
g120 and 463(88) ; 3017(169)
g121 and 463(88) 456(94) ; 621(170)
g122 and 3087(90) ; 3093(171)
g123 and 3079(91) ; 3085(172)
g124 and 456(94) ; 3010(173)
g125 and 3007(97) ; 3013(174)
g126 and 442(98) ; 636(175)
g127 and 45(5) 732(117) 717(120) ; 896(176)
g128 and 802(100) ; 657(177)
g129 and 802(100) ; 675(178)
g130 and 791(103) 799(101) 714(124) ; 816(179)
g131 and 799(101) 704(126) ; 823(180)
g132 and 798(102) 714(124) ; 807(181)
g133 and 791(103) ; 794(182)
g134 and 1699(105) ; 1717(183)
g135 and 1699(105) ; 1724(184)
g136 and 1699(105) ; 1731(185)
g137 and 1699(105) ; 1738(186)
g138 and 1699(105) ; 1745(187)
g139 and 1699(105) ; 1752(188)
g140 and 1699(105) ; 1759(189)
g141 and 1699(105) ; 1766(190)
g142 and 780(106) ; 784(191)
g143 and 780(106) ; 1681(192)
g144 and 776(107) ; 1512(193)
g145 and 788(109) ; 1790(194)
g146 and 788(109) ; 1808(195)
g147 and 1051(112) ; 1054(196)
g148 and 1051(112) ; 1057(197)
g149 and 20(2)* 758(108)* ; 759(198)
g150 and 741(116) ; 973(199)
g151 and 741(116) ; 980(200)
g152 and 741(116) ; 987(201)
g153 and 741(116) ; 994(202)
g154 and 741(116) ; 1001(203)
g155 and 741(116) ; 1008(204)
g156 and 741(116) ; 1015(205)
g157 and 741(116) ; 1022(206)
g158 and 732(117) 717(120) 704(126) ; 2278(207)
g159 and 736(118) 724(119) 707(127) ; 860(208)
g160 and 736(118) 724(119) 707(127) ; 861(209)
g161 and 724(119) 707(127) ; 864(210)
g162 and 717(120) ; 721(211)
g163 and 731(121) ; 1772(212)
g164 and 1(0)* 2051(104)* ; 2052(213)
g165 and 1(0)* 1828(110)* ; 1829(214)
g166 and 1827(122) 1826(123) ; 1834(215)
g167 and 890(125) ; 893(216)
g168 and 2874(129) ; 2877(217)
g169 and 2963(133) 2960(52) ; 2965(218)
g170 and 552(132) 551(134) 550(136) 549(139) ; 554(219)
g171 and 2964(131) 2957(53) ; 2966(220)
g172 and 1766(190) 257(34) ; 1769(221)
g173 and 2953(138) 2950(55) ; 2955(222)
g174 and 1759(189) 250(33) ; 1762(223)
g175 and 2954(135) 2947(56) ; 2956(224)
g176 and 1752(188) 244(32) ; 1755(225)
g177 and 2945(142) 2942(57) ; 560(226)
g178 and 548(141) 547(143) 546(145) 545(147) ; 553(227)
g179 and 1745(187) 238(31) ; 1748(228)
g180 and 2946(140) 2939(58) ; 561(229)
g181 and 1738(186) 232(30) ; 1741(230)
g182 and 2937(146) 2934(59) ; 555(231)
g183 and 1731(185) 226(29) ; 1734(232)
g184 and 2938(144) 2931(60) ; 556(233)
g185 and 1724(184) 223(28) ; 1727(234)
g186 and 1717(183) 222(27) ; 1720(235)
g187 and 343(47) 213(26) 2278(207) ; 2302(236)
g188 and 343(47) 213(26) 2278(207) ; 2298(237)
g189 and 343(47) 213(26) 2278(207) ; 2293(238)
g190 and 343(47) 213(26) 2278(207) ; 2289(239)
g191 and 213(26) 2278(207) ; 2288(240)
g192 and 213(26) 2278(207) ; 2285(241)
g193 and 1054(196) 1048(62) ; 1063(242)
g194 and 1054(196) 200(25) ; 1060(243)
g195 and 1022(206) 116(13) ; 1025(244)
g196 and 3040(152) ; 3044(245)
g197 and 905(155) 540(65) ; 630(246)
g198 and 905(155) 540(65) ; 634(247)
g199 and 3101(160) 3098(153) ; 646(248)
g200 and 3098(153) ; 3102(249)
g201 and 3109(159) 3106(154) ; 912(250)
g202 and 3106(154) ; 3110(251)
g203 and 1001(203) 906(156) ; 1004(252)
g204 and 1015(205) 851(68) ; 1018(253)
g205 and 3037(157) ; 3043(254)
g206 and 3030(161) ; 3034(255)
g207 and 626(158) 87(10) ; 654(256)
g208 and 626(158) 87(10) ; 354(257)
g209 and 3027(162) ; 3033(258)
g210 and 994(202) 77(9) ; 997(259)
g211 and 625(167) 479(82) ; 352(260)
g212 and 3020(163) ; 3024(261)
g213 and 3085(172) 3082(165) ; 642(262)
g214 and 3082(165) ; 3086(263)
g215 and 3093(171) 3090(166) ; 903(264)
g216 and 3090(166) ; 3094(265)
g217 and 973(199) 897(168) ; 976(266)
g218 and 987(201) 836(85) ; 990(267)
g219 and 3017(169) ; 3023(268)
g220 and 636(175) 460(89) ; 644(269)
g221 and 3013(174) 3010(173) ; 3015(270)
g222 and 3010(173) ; 3014(271)
g223 and 636(175) ; 639(272)
g224 and 621(170) 432(99) ; 650(273)
g225 and 657(177) ; 660(274)
g226 and 675(178) ; 678(275)
g227 and 816(179) ; 2128(276)
g228 and 816(179) ; 2181(277)
g229 and 816(179) ; 2233(278)
g230 and 823(180) ; 2076(279)
g231 and 807(181) ; 1870(280)
g232 and 807(181) ; 1920(281)
g233 and 807(181) ; 1971(282)
g234 and 807(181) ; 2021(283)
g235 and 794(182) 784(191) ; 1527(284)
g236 and 1699(105) 1681(192) ; 1718(285)
g237 and 1699(105) 1681(192) ; 1725(286)
g238 and 1699(105) 1681(192) ; 1732(287)
g239 and 1699(105) 1681(192) ; 1739(288)
g240 and 1699(105) 1681(192) ; 1746(289)
g241 and 1699(105) 1681(192) ; 1753(290)
g242 and 1699(105) 1681(192) ; 1760(291)
g243 and 1699(105) 1681(192) ; 1767(292)
g244 and 780(106) 860(208) ; 806(293)
g245 and 1681(192) ; 1716(294)
g246 and 1681(192) ; 1723(295)
g247 and 1681(192) ; 1730(296)
g248 and 1681(192) ; 1737(297)
g249 and 1681(192) ; 1744(298)
g250 and 1681(192) ; 1751(299)
g251 and 1681(192) ; 1758(300)
g252 and 1681(192) ; 1765(301)
g253 and 794(182) 776(107) ; 1530(302)
g254 and 776(107) 860(208) ; 804(303)
g255 and 1512(193) ; 1581(304)
g256 and 1512(193) ; 1585(305)
g257 and 1512(193) ; 1589(306)
g258 and 1512(193) ; 1593(307)
g259 and 1512(193) ; 1597(308)
g260 and 1512(193) ; 1601(309)
g261 and 1512(193) ; 1605(310)
g262 and 1057(197) 1050(113) ; 1069(311)
g263 and 1057(197) 1049(114) ; 1066(312)
g264 and 759(198) ; 974(313)
g265 and 759(198) ; 981(314)
g266 and 759(198) ; 988(315)
g267 and 759(198) ; 995(316)
g268 and 759(198) ; 1002(317)
g269 and 759(198) ; 1009(318)
g270 and 759(198) ; 1016(319)
g271 and 759(198) ; 1023(320)
g272 and 759(198) 741(116) ; 975(321)
g273 and 759(198) 741(116) ; 982(322)
g274 and 759(198) 741(116) ; 989(323)
g275 and 759(198) 741(116) ; 996(324)
g276 and 759(198) 741(116) ; 1003(325)
g277 and 759(198) 741(116) ; 1010(326)
g278 and 759(198) 741(116) ; 1017(327)
g279 and 759(198) 741(116) ; 1024(328)
g280 and 784(191) 732(117) 724(119) ; 1563(329)
g281 and 736(118) 721(211) 707(127) ; 855(330)
g282 and 861(209) ; 915(331)
g283 and 794(182) 736(118) 724(119) 707(127) ; 867(332)
g284 and 864(210) ; 941(333)
g285 and 784(191) 724(119) ; 1572(334)
g286 and 1834(215) ; 1851(335)
g287 and 1834(215) ; 1901(336)
g288 and 1834(215) ; 1952(337)
g289 and 1834(215) ; 2002(338)
g290 and 1834(215) ; 2057(339)
g291 and 1834(215) ; 2109(340)
g292 and 1834(215) ; 2162(341)
g293 and 1834(215) ; 2214(342)
g294 and 1808(195) 13(1) 1(0) ; 1809(343)
g295 and 1790(194) 13(1) 1(0) ; 1791(344)
g296 and 1772(212)* 1(0)* ; 1773(345)
g297 and 896(176) 890(125) ; 956(346)
g298 and 893(216) ; 927(347)
g299 and 1541(151) 721(211) 707(127) ; 1542(348)
g300 and 2897(49) 2877(217) ; 2903(349)
g301 and 2897(49) 2877(217) ; 2900(350)
g302 and 1765(301) 303(40) ; 1768(351)
g303 and 1758(300) 294(39) ; 1761(352)
g304 and 1751(299) 283(38) ; 1754(353)
g305 and 1023(320) 283(38) ; 1026(354)
g306 and 2966(220) 2965(218) ; 2986(355)
g307 and 554(219) 553(227) ; 586(356)
g308 and 1767(292) 264(35) ; 1770(357)
g309 and 1760(291) 257(34) ; 1763(358)
g310 and 2956(224) 2955(222) ; 2983(359)
g311 and 1753(290) 250(33) ; 1756(360)
g312 and 915(331) 588(137) ; 920(361)
g313 and 1746(289) 244(32) ; 1749(362)
g314 and 561(229) 560(226) ; 562(363)
g315 and 1739(288) 238(31) ; 1742(364)
g316 and 1732(287) 232(30) ; 1735(365)
g317 and 556(233) 555(231) ; 557(366)
g318 and 1725(286) 226(29) ; 1728(367)
g319 and 1718(285) 223(28) ; 1721(368)
g320 and 2293(238) ; 2485(369)
g321 and 1069(311) 1038(148) ; 1096(370)
g322 and 1066(312) 1038(148) ; 1108(371)
g323 and 1063(242) 1038(148) ; 1144(372)
g324 and 1060(243) 1038(148) ; 1156(373)
g325 and 1069(311) 1043(149) ; 1072(374)
g326 and 1066(312) 1043(149) ; 1084(375)
g327 and 1063(242) 1043(149) ; 1120(376)
g328 and 1060(243) 1043(149) ; 1132(377)
g329 and 982(322) 159(21) ; 985(378)
g330 and 975(321) 150(20) ; 978(379)
g331 and 1773(345)* 116(13)* ; 2219(380)
g332 and 1744(298) 116(13) ; 1747(381)
g333 and 1016(319) 116(13) ; 1019(382)
g334 and 3043(254) 3040(152) ; 3045(383)
g335 and 1773(345)* 107(12)* ; 2167(384)
g336 and 1737(297) 107(12) ; 1740(385)
g337 and 1009(318) 107(12) ; 1012(386)
g338 and 3044(245) 3037(157) ; 3046(387)
g339 and 1773(345)* 97(11)* ; 2114(388)
g340 and 1730(296) 97(11) ; 1733(389)
g341 and 3110(251) 3103(71) ; 913(390)
g342 and 3102(249) 3095(72) ; 647(391)
g343 and 1002(317) 845(74) ; 1005(392)
g344 and 1024(328) 845(74) ; 1027(393)
g345 and 3033(258) 3030(161) ; 3035(394)
g346 and 1773(345)* 87(10)* ; 2062(395)
g347 and 1723(295) 87(10) ; 1726(396)
g348 and 995(316) 839(78) ; 998(397)
g349 and 1017(327) 839(78) ; 1020(398)
g350 and 354(257) ; 355(399)
g351 and 3034(255) 3027(162) ; 3036(400)
g352 and 1773(345)* 77(9)* ; 2007(401)
g353 and 1716(294) 77(9) ; 1719(402)
g354 and 1010(326) 77(9) ; 1013(403)
g355 and 988(315) 77(9) ; 991(404)
g356 and 352(260) ; 353(405)
g357 and 3023(268) 3020(163) ; 3025(406)
g358 and 1773(345)* 68(8)* ; 1957(407)
g359 and 981(314) 833(86) ; 984(408)
g360 and 1003(325) 833(86) ; 1006(409)
g361 and 3024(261) 3017(169) ; 3026(410)
g362 and 1773(345)* 58(7)* ; 1906(411)
g363 and 3094(265) 3087(90) ; 904(412)
g364 and 3086(263) 3079(91) ; 643(413)
g365 and 974(313) 828(93) ; 977(414)
g366 and 996(324) 828(93) ; 999(415)
g367 and 58(7) 442(98) 635(164) 630(246) ; 655(416)
g368 and 1773(345)* 50(6)* ; 1856(417)
g369 and 989(323) 50(6) ; 992(418)
g370 and 3014(271) 3007(97) ; 3016(419)
g371 and 675(178) 650(273) ; 680(420)
g372 and 1527(284) ; 1533(421)
g373 and 1530(302) 1527(284) ; 1535(422)
g374 and 806(293) 804(303) ; 613(423)
g375 and 806(293) ; 616(424)
g376 and 806(293) 804(303) ; 668(425)
g377 and 806(293) ; 671(426)
g378 and 806(293) ; 685(427)
g379 and 806(293) 804(303) ; 688(428)
g380 and 806(293) ; 696(429)
g381 and 806(293) 804(303) ; 699(430)
g382 and 1530(302) ; 1534(431)
g383 and 804(303) ; 610(432)
g384 and 804(303) ; 665(433)
g385 and 804(303) ; 683(434)
g386 and 804(303) ; 694(435)
g387 and 1563(329) ; 1646(436)
g388 and 1563(329) ; 1655(437)
g389 and 1563(329) ; 1664(438)
g390 and 1563(329) ; 1673(439)
g391 and 855(330) ; 914(440)
g392 and 855(330) ; 942(441)
g393 and 861(209) 855(330) ; 916(442)
g394 and 867(332) ; 870(443)
g395 and 867(332) ; 887(444)
g396 and 855(330) 864(210) ; 943(445)
g397 and 1572(334) ; 1610(446)
g398 and 1572(334) ; 1619(447)
g399 and 1572(334) ; 1628(448)
g400 and 1572(334) ; 1637(449)
g401 and 1773(345) 1834(215) ; 1852(450)
g402 and 1773(345) 1834(215) ; 1902(451)
g403 and 1773(345) 1834(215) ; 1953(452)
g404 and 1773(345) 1834(215) ; 2003(453)
g405 and 1773(345) 1834(215) ; 2058(454)
g406 and 1773(345) 1834(215) ; 2110(455)
g407 and 1773(345) 1834(215) ; 2163(456)
g408 and 1773(345) 1834(215) ; 2215(457)
g409 and 1809(343) ; 1812(458)
g410 and 1809(343) ; 1817(459)
g411 and 1791(344) ; 1794(460)
g412 and 1791(344) ; 1799(461)
g413 and 956(346) ; 2678(462)
g414 and 956(346) ; 2697(463)
g415 and 956(346) ; 2716(464)
g416 and 956(346) ; 2733(465)
g417 and 956(346) ; 2751(466)
g418 and 956(346) ; 2768(467)
g419 and 956(346) ; 2785(468)
g420 and 956(346) ; 2802(469)
g421 and 1542(348) ; 1545(470)
g422 and 1542(348) ; 1554(471)
g423 and 816(179) 274(37) 1799(461) ; 2235(472)
g424 and 816(179) 274(37) 1799(461) ; 2183(473)
g425 and 816(179) 274(37) 1799(461) ; 2130(474)
g426 and 823(180) 274(37) 1799(461) ; 2078(475)
g427 and 807(181) 274(37) 1817(459) ; 2023(476)
g428 and 807(181) 274(37) 1817(459) ; 1973(477)
g429 and 807(181) 274(37) 1817(459) ; 1922(478)
g430 and 807(181) 274(37) 1817(459) ; 1872(479)
g431 and 2233(278) 270(36) 1799(461) ; 2234(480)
g432 and 2986(355) ; 2990(481)
g433 and 916(442) 586(356) ; 923(482)
g434 and 2181(277) 264(35) 1799(461) ; 2182(483)
g435 and 2128(276) 257(34) 1799(461) ; 2129(484)
g436 and 1770(357)* 1769(221)* 1768(351)* ; 1771(485)
g437 and 2983(359) ; 2989(486)
g438 and 2076(279) 250(33) 1799(461) ; 2077(487)
g439 and 1763(358)* 1762(223)* 1761(352)* ; 1764(488)
g440 and 2021(283) 244(32) 1817(459) ; 2022(489)
g441 and 1756(360)* 1755(225)* 1754(353)* ; 1757(490)
g442 and 562(363) ; 2970(491)
g443 and 562(363) ; 2978(492)
g444 and 1971(282) 238(31) 1817(459) ; 1972(493)
g445 and 1749(362)* 1748(228)* 1747(381)* ; 1750(494)
g446 and 1920(281) 232(30) 1817(459) ; 1921(495)
g447 and 1742(364)* 1741(230)* 1740(385)* ; 1743(496)
g448 and 557(366) ; 2967(497)
g449 and 557(366) ; 2975(498)
g450 and 1870(280) 226(29) 1817(459) ; 1871(499)
g451 and 1735(365)* 1734(232)* 1733(389)* ; 1736(500)
g452 and 1728(367)* 1727(234)* 1726(396)* ; 1729(501)
g453 and 1721(368)* 1720(235)* 1719(402)* ; 1722(502)
g454 and 2485(369) ; 2488(503)
g455 and 1096(370) ; 1099(504)
g456 and 1096(370) ; 1186(505)
g457 and 1108(371) ; 1111(506)
g458 and 1108(371) ; 1195(507)
g459 and 1144(372) ; 1147(508)
g460 and 1144(372) ; 1222(509)
g461 and 1156(373) ; 1159(510)
g462 and 1156(373) ; 1231(511)
g463 and 1072(374) ; 1075(512)
g464 and 1072(374) ; 1168(513)
g465 and 1084(375) ; 1087(514)
g466 and 1084(375) ; 1177(515)
g467 and 1120(376) ; 1123(516)
g468 and 1120(376) ; 1204(517)
g469 and 1132(377) ; 1135(518)
g470 and 1132(377) ; 1213(519)
g471 and 2215(457) 2052(213) 116(13) ; 2222(520)
g472 and 1027(393)* 1026(354)* 1025(244)* ; 1028(521)
g473 and 3046(387) 3045(383) ; 3058(522)
g474 and 696(429) 634(247) ; 701(523)
g475 and 688(428) 540(65) ; 691(524)
g476 and 2163(456) 2052(213) 107(12) ; 2170(525)
g477 and 647(391) 646(248) ; 648(526)
g478 and 913(390) 912(250) ; 910(527)
g479 and 1006(409)* 1005(392)* 1004(252)* ; 1007(528)
g480 and 1020(398)* 1019(382)* 1018(253)* ; 1021(529)
g481 and 699(430) 526(69) ; 702(530)
g482 and 2110(455) 2052(213) 97(11) ; 2117(531)
g483 and 3036(400) 3035(394) ; 3055(532)
g484 and 668(425) 513(75) ; 672(533)
g485 and 2058(454) 2052(213) 87(10) ; 2065(534)
g486 and 685(427) 654(256) ; 690(535)
g487 and 613(423) 501(79) ; 617(536)
g488 and 2003(453) 1829(214) 77(9) ; 2010(537)
g489 and 999(415)* 998(397)* 997(259)* ; 1000(538)
g490 and 3026(410) 3025(406) ; 3050(539)
g491 and 1953(452) 1829(214) 68(8) ; 1960(540)
g492 and 643(413) 642(262) ; 640(541)
g493 and 904(412) 903(264) ; 901(542)
g494 and 978(379)* 977(414)* 976(266)* ; 979(543)
g495 and 992(418)* 991(404)* 990(267)* ; 993(544)
g496 and 1902(451) 1829(214) 58(7) ; 1909(545)
g497 and 3016(419) 3015(270) ; 3047(546)
g498 and 1852(450) 1829(214) 50(6) ; 1859(547)
g499 and 1535(422) 442(98) ; 1538(548)
g500 and 914(440) 650(273) ; 917(549)
g501 and 657(177) 655(416) ; 662(550)
g502 and 1563(329) 1554(471) ; 1647(551)
g503 and 1563(329) 1554(471) ; 1656(552)
g504 and 1563(329) 1554(471) ; 1665(553)
g505 and 1563(329) 1554(471) ; 1674(554)
g506 and 870(443) ; 2679(555)
g507 and 870(443) ; 2698(556)
g508 and 870(443) ; 2717(557)
g509 and 870(443) ; 2734(558)
g510 and 870(443) ; 2752(559)
g511 and 870(443) ; 2769(560)
g512 and 870(443) ; 2786(561)
g513 and 870(443) ; 2803(562)
g514 and 887(444) ; 926(563)
g515 and 1572(334) 1545(470) ; 1611(564)
g516 and 1572(334) 1545(470) ; 1620(565)
g517 and 1572(334) 1545(470) ; 1629(566)
g518 and 1572(334) 1545(470) ; 1638(567)
g519 and 870(443) 956(346) ; 2680(568)
g520 and 870(443) 956(346) ; 2699(569)
g521 and 870(443) 956(346) ; 2718(570)
g522 and 870(443) 956(346) ; 2735(571)
g523 and 870(443) 956(346) ; 2753(572)
g524 and 870(443) 956(346) ; 2770(573)
g525 and 870(443) 956(346) ; 2787(574)
g526 and 870(443) 956(346) ; 2804(575)
g527 and 893(216) 887(444) ; 928(576)
g528 and 1545(470) ; 1609(577)
g529 and 1545(470) ; 1618(578)
g530 and 1545(470) ; 1627(579)
g531 and 1545(470) ; 1636(580)
g532 and 1554(471) ; 1645(581)
g533 and 1554(471) ; 1654(582)
g534 and 1554(471) ; 1663(583)
g535 and 1554(471) ; 1672(584)
g536 and 2989(486) 2986(355) ; 574(585)
g537 and 2990(481) 2983(359) ; 575(586)
g538 and 923(482)* 920(361)* 917(549)* ; 359(587)
g539 and 923(482)* 920(361)* 917(549)* ; 1029(588)
g540 and 2970(491) ; 2974(589)
g541 and 2978(492) ; 2982(590)
g542 and 2967(497) ; 2973(591)
g543 and 2975(498) ; 2981(592)
g544 and 1099(504) ; 1242(593)
g545 and 1099(504) ; 1259(594)
g546 and 1099(504) ; 1276(595)
g547 and 1099(504) ; 1293(596)
g548 and 1099(504) ; 1310(597)
g549 and 1099(504) ; 1327(598)
g550 and 1099(504) ; 1344(599)
g551 and 1099(504) ; 1361(600)
g552 and 1186(505) ; 1378(601)
g553 and 1186(505) ; 1395(602)
g554 and 1186(505) ; 1412(603)
g555 and 1186(505) ; 1429(604)
g556 and 1186(505) ; 1446(605)
g557 and 1186(505) ; 1463(606)
g558 and 1186(505) ; 1480(607)
g559 and 1186(505) ; 1497(608)
g560 and 1111(506) ; 1243(609)
g561 and 1111(506) ; 1260(610)
g562 and 1111(506) ; 1277(611)
g563 and 1111(506) ; 1294(612)
g564 and 1111(506) ; 1311(613)
g565 and 1111(506) ; 1328(614)
g566 and 1111(506) ; 1345(615)
g567 and 1111(506) ; 1362(616)
g568 and 1195(507) ; 1379(617)
g569 and 1195(507) ; 1396(618)
g570 and 1195(507) ; 1413(619)
g571 and 1195(507) ; 1430(620)
g572 and 1195(507) ; 1447(621)
g573 and 1195(507) ; 1464(622)
g574 and 1195(507) ; 1481(623)
g575 and 1195(507) ; 1498(624)
g576 and 1147(508) ; 1246(625)
g577 and 1147(508) ; 1263(626)
g578 and 1147(508) ; 1280(627)
g579 and 1147(508) ; 1297(628)
g580 and 1147(508) ; 1314(629)
g581 and 1147(508) ; 1331(630)
g582 and 1147(508) ; 1348(631)
g583 and 1147(508) ; 1365(632)
g584 and 1222(509) ; 1382(633)
g585 and 1222(509) ; 1399(634)
g586 and 1222(509) ; 1416(635)
g587 and 1222(509) ; 1433(636)
g588 and 1222(509) ; 1450(637)
g589 and 1222(509) ; 1467(638)
g590 and 1222(509) ; 1484(639)
g591 and 1222(509) ; 1501(640)
g592 and 1159(510) ; 1247(641)
g593 and 1159(510) ; 1264(642)
g594 and 1159(510) ; 1281(643)
g595 and 1159(510) ; 1298(644)
g596 and 1159(510) ; 1315(645)
g597 and 1159(510) ; 1332(646)
g598 and 1159(510) ; 1349(647)
g599 and 1159(510) ; 1366(648)
g600 and 1231(511) ; 1383(649)
g601 and 1231(511) ; 1400(650)
g602 and 1231(511) ; 1417(651)
g603 and 1231(511) ; 1434(652)
g604 and 1231(511) ; 1451(653)
g605 and 1231(511) ; 1468(654)
g606 and 1231(511) ; 1485(655)
g607 and 1231(511) ; 1502(656)
g608 and 1075(512) ; 1240(657)
g609 and 1075(512) ; 1257(658)
g610 and 1075(512) ; 1274(659)
g611 and 1075(512) ; 1291(660)
g612 and 1075(512) ; 1308(661)
g613 and 1075(512) ; 1325(662)
g614 and 1075(512) ; 1342(663)
g615 and 1075(512) ; 1359(664)
g616 and 1168(513) ; 1376(665)
g617 and 1168(513) ; 1393(666)
g618 and 1168(513) ; 1410(667)
g619 and 1168(513) ; 1427(668)
g620 and 1168(513) ; 1444(669)
g621 and 1168(513) ; 1461(670)
g622 and 1168(513) ; 1478(671)
g623 and 1168(513) ; 1495(672)
g624 and 1087(514) ; 1241(673)
g625 and 1087(514) ; 1258(674)
g626 and 1087(514) ; 1275(675)
g627 and 1087(514) ; 1292(676)
g628 and 1087(514) ; 1309(677)
g629 and 1087(514) ; 1326(678)
g630 and 1087(514) ; 1343(679)
g631 and 1087(514) ; 1360(680)
g632 and 1177(515) ; 1377(681)
g633 and 1177(515) ; 1394(682)
g634 and 1177(515) ; 1411(683)
g635 and 1177(515) ; 1428(684)
g636 and 1177(515) ; 1445(685)
g637 and 1177(515) ; 1462(686)
g638 and 1177(515) ; 1479(687)
g639 and 1177(515) ; 1496(688)
g640 and 1123(516) ; 1244(689)
g641 and 1123(516) ; 1261(690)
g642 and 1123(516) ; 1278(691)
g643 and 1123(516) ; 1295(692)
g644 and 1123(516) ; 1312(693)
g645 and 1123(516) ; 1329(694)
g646 and 1123(516) ; 1346(695)
g647 and 1123(516) ; 1363(696)
g648 and 1204(517) ; 1380(697)
g649 and 1204(517) ; 1397(698)
g650 and 1204(517) ; 1414(699)
g651 and 1204(517) ; 1431(700)
g652 and 1204(517) ; 1448(701)
g653 and 1204(517) ; 1465(702)
g654 and 1204(517) ; 1482(703)
g655 and 1204(517) ; 1499(704)
g656 and 1135(518) ; 1245(705)
g657 and 1135(518) ; 1262(706)
g658 and 1135(518) ; 1279(707)
g659 and 1135(518) ; 1296(708)
g660 and 1135(518) ; 1313(709)
g661 and 1135(518) ; 1330(710)
g662 and 1135(518) ; 1347(711)
g663 and 1135(518) ; 1364(712)
g664 and 1213(519) ; 1381(713)
g665 and 1213(519) ; 1398(714)
g666 and 1213(519) ; 1415(715)
g667 and 1213(519) ; 1432(716)
g668 and 1213(519) ; 1449(717)
g669 and 1213(519) ; 1466(718)
g670 and 1213(519) ; 1483(719)
g671 and 1213(519) ; 1500(720)
g672 and 3058(522) ; 3062(721)
g673 and 928(576) 630(246) ; 938(722)
g674 and 648(526) 530(66) ; 649(723)
g675 and 910(527) ; 911(724)
g676 and 3055(532) ; 3061(725)
g677 and 3050(539) ; 3054(726)
g678 and 1638(567) 479(82) ; 1643(727)
g679 and 639(272) 476(83) 640(541) ; 641(728)
g680 and 901(542) ; 902(729)
g681 and 1629(566) 463(88) ; 1634(730)
g682 and 3047(546) ; 3053(731)
g683 and 1620(565) 456(94) ; 1625(732)
g684 and 1611(564) 442(98) ; 1616(733)
g685 and 926(563) 650(273) ; 929(734)
g686 and 1851(335) 979(543) ; 1853(735)
g687 and 1952(337) 993(544) ; 1954(736)
g688 and 2002(338) 1000(538) ; 2004(737)
g689 and 2057(339) 1007(528) ; 2059(738)
g690 and 2162(341) 1021(529) ; 2164(739)
g691 and 2214(342) 1028(521) ; 2216(740)
g692 and 1722(502) 1812(458) ; 1873(741)
g693 and 1729(501) 1812(458) ; 1923(742)
g694 and 1736(500) 1812(458) ; 1974(743)
g695 and 1743(496) 1812(458) ; 2024(744)
g696 and 1750(494) 1794(460) ; 2079(745)
g697 and 1757(490) 1794(460) ; 2131(746)
g698 and 1764(488) 1794(460) ; 2184(747)
g699 and 1771(485) 1794(460) ; 2236(748)
g700 and 1495(672) 329(45) ; 1503(749)
g701 and 1502(656) 326(44) ; 1510(750)
g702 and 1478(671) 326(44) ; 1486(751)
g703 and 1501(640) 322(43) ; 1509(752)
g704 and 1485(655) 322(43) ; 1493(753)
g705 and 1461(670) 322(43) ; 1469(754)
g706 and 1500(720) 317(42) ; 1508(755)
g707 and 1484(639) 317(42) ; 1492(756)
g708 and 1468(654) 317(42) ; 1476(757)
g709 and 1444(669) 317(42) ; 1452(758)
g710 and 1499(704) 311(41) ; 1507(759)
g711 and 1483(719) 311(41) ; 1491(760)
g712 and 1467(638) 311(41) ; 1475(761)
g713 and 1451(653) 311(41) ; 1459(762)
g714 and 1427(668) 311(41) ; 1435(763)
g715 and 1498(624) 303(40) ; 1506(764)
g716 and 1482(703) 303(40) ; 1490(765)
g717 and 1466(718) 303(40) ; 1474(766)
g718 and 1450(637) 303(40) ; 1458(767)
g719 and 1434(652) 303(40) ; 1442(768)
g720 and 1410(667) 303(40) ; 1418(769)
g721 and 1497(608) 294(39) ; 1505(770)
g722 and 1481(623) 294(39) ; 1489(771)
g723 and 1465(702) 294(39) ; 1473(772)
g724 and 1449(717) 294(39) ; 1457(773)
g725 and 1433(636) 294(39) ; 1441(774)
g726 and 1417(651) 294(39) ; 1425(775)
g727 and 1393(666) 294(39) ; 1401(776)
g728 and 1496(688) 283(38) ; 1504(777)
g729 and 1480(607) 283(38) ; 1488(778)
g730 and 1464(622) 283(38) ; 1472(779)
g731 and 1448(701) 283(38) ; 1456(780)
g732 and 1432(716) 283(38) ; 1440(781)
g733 and 1416(635) 283(38) ; 1424(782)
g734 and 1400(650) 283(38) ; 1408(783)
g735 and 1376(665) 283(38) ; 1384(784)
g736 and 2236(748)* 2235(472)* 2234(480)* ; 2237(785)
g737 and 2184(747)* 2183(473)* 2182(483)* ; 2185(786)
g738 and 2131(746)* 2130(474)* 2129(484)* ; 2132(787)
g739 and 2079(745)* 2078(475)* 2077(487)* ; 2080(788)
g740 and 2024(744)* 2023(476)* 2022(489)* ; 2025(789)
g741 and 1974(743)* 1973(477)* 1972(493)* ; 1975(790)
g742 and 1923(742)* 1922(478)* 1921(495)* ; 1924(791)
g743 and 1873(741)* 1872(479)* 1871(499)* ; 1874(792)
g744 and 575(586) 574(585) ; 576(793)
g745 and 1029(588) ; 360(794)
g746 and 2973(591) 2970(491) ; 565(795)
g747 and 2981(592) 2978(492) ; 569(796)
g748 and 2974(589) 2967(497) ; 566(797)
g749 and 2982(590) 2975(498) ; 570(798)
g750 and 1359(664) 159(21) ; 1367(799)
g751 and 1349(647) 159(21) ; 1357(800)
g752 and 1331(630) 159(21) ; 1339(801)
g753 and 1313(709) 159(21) ; 1321(802)
g754 and 1295(692) 159(21) ; 1303(803)
g755 and 1277(611) 159(21) ; 1285(804)
g756 and 1259(594) 159(21) ; 1267(805)
g757 and 1241(673) 159(21) ; 1249(806)
g758 and 1342(663) 150(20) ; 1350(807)
g759 and 1332(646) 150(20) ; 1340(808)
g760 and 1314(629) 150(20) ; 1322(809)
g761 and 1296(708) 150(20) ; 1304(810)
g762 and 1278(691) 150(20) ; 1286(811)
g763 and 1260(610) 150(20) ; 1268(812)
g764 and 1242(593) 150(20) ; 1250(813)
g765 and 1325(662) 143(19) ; 1333(814)
g766 and 1315(645) 143(19) ; 1323(815)
g767 and 1297(628) 143(19) ; 1305(816)
g768 and 1279(707) 143(19) ; 1287(817)
g769 and 1261(690) 143(19) ; 1269(818)
g770 and 1243(609) 143(19) ; 1251(819)
g771 and 1308(661) 137(18) ; 1316(820)
g772 and 1298(644) 137(18) ; 1306(821)
g773 and 1280(627) 137(18) ; 1288(822)
g774 and 1262(706) 137(18) ; 1270(823)
g775 and 1244(689) 137(18) ; 1252(824)
g776 and 1291(660) 132(17) ; 1299(825)
g777 and 1281(643) 132(17) ; 1289(826)
g778 and 1263(626) 132(17) ; 1271(827)
g779 and 1245(705) 132(17) ; 1253(828)
g780 and 1274(659) 128(16) ; 1282(829)
g781 and 1264(642) 128(16) ; 1272(830)
g782 and 1246(625) 128(16) ; 1254(831)
g783 and 1257(658) 125(15) ; 1265(832)
g784 and 1247(641) 125(15) ; 1255(833)
g785 and 1240(657) 124(14) ; 1248(834)
g786 and 2222(520)* 2219(380)* 2216(740)* ; 2225(835)
g787 and 2222(520)* 2219(380)* 2216(740)* ; 2229(836)
g788 and 3061(725) 3058(522) ; 595(837)
g789 and 1383(649) 530(66) ; 1391(838)
g790 and 1399(634) 530(66) ; 1407(839)
g791 and 1415(715) 530(66) ; 1423(840)
g792 and 1431(700) 530(66) ; 1439(841)
g793 and 1447(621) 530(66) ; 1455(842)
g794 and 1463(606) 530(66) ; 1471(843)
g795 and 1479(687) 530(66) ; 1487(844)
g796 and 2170(525)* 2167(384)* 2164(739)* ; 2173(845)
g797 and 2170(525)* 2167(384)* 2164(739)* ; 2177(846)
g798 and 1360(680) 517(70) ; 1368(847)
g799 and 1382(633) 517(70) ; 1390(848)
g800 and 1398(714) 517(70) ; 1406(849)
g801 and 1414(699) 517(70) ; 1422(850)
g802 and 1430(620) 517(70) ; 1438(851)
g803 and 1446(605) 517(70) ; 1454(852)
g804 and 1462(686) 517(70) ; 1470(853)
g805 and 3062(721) 3055(532) ; 596(854)
g806 and 1343(679) 504(76) ; 1351(855)
g807 and 1361(600) 504(76) ; 1369(856)
g808 and 1381(713) 504(76) ; 1389(857)
g809 and 1397(698) 504(76) ; 1405(858)
g810 and 1413(619) 504(76) ; 1421(859)
g811 and 1429(604) 504(76) ; 1437(860)
g812 and 1445(685) 504(76) ; 1453(861)
g813 and 2065(534)* 2062(395)* 2059(738)* ; 2068(862)
g814 and 2065(534)* 2062(395)* 2059(738)* ; 2072(863)
g815 and 1326(678) 492(80) ; 1334(864)
g816 and 1344(599) 492(80) ; 1352(865)
g817 and 1362(616) 492(80) ; 1370(866)
g818 and 1380(697) 492(80) ; 1388(867)
g819 and 1396(618) 492(80) ; 1404(868)
g820 and 1412(603) 492(80) ; 1420(869)
g821 and 1428(684) 492(80) ; 1436(870)
g822 and 2010(537)* 2007(401)* 2004(737)* ; 2013(871)
g823 and 2010(537)* 2007(401)* 2004(737)* ; 2017(872)
g824 and 1309(677) 483(81) ; 1317(873)
g825 and 1327(598) 483(81) ; 1335(874)
g826 and 1345(615) 483(81) ; 1353(875)
g827 and 1363(696) 483(81) ; 1371(876)
g828 and 1379(617) 483(81) ; 1387(877)
g829 and 1395(602) 483(81) ; 1403(878)
g830 and 1411(683) 483(81) ; 1419(879)
g831 and 3053(731) 3050(539) ; 589(880)
g832 and 1960(540)* 1957(407)* 1954(736)* ; 1963(881)
g833 and 1960(540)* 1957(407)* 1954(736)* ; 1967(882)
g834 and 1292(676) 467(87) ; 1300(883)
g835 and 1310(597) 467(87) ; 1318(884)
g836 and 1328(614) 467(87) ; 1336(885)
g837 and 1346(695) 467(87) ; 1354(886)
g838 and 1364(712) 467(87) ; 1372(887)
g839 and 1378(601) 467(87) ; 1386(888)
g840 and 1394(682) 467(87) ; 1402(889)
g841 and 644(269)* 641(728)* ; 645(890)
g842 and 3054(726) 3047(546) ; 590(891)
g843 and 1275(675) 447(95) ; 1283(892)
g844 and 1293(596) 447(95) ; 1301(893)
g845 and 1311(613) 447(95) ; 1319(894)
g846 and 1329(694) 447(95) ; 1337(895)
g847 and 1347(711) 447(95) ; 1355(896)
g848 and 1365(632) 447(95) ; 1373(897)
g849 and 1377(681) 447(95) ; 1385(898)
g850 and 1859(547)* 1856(417)* 1853(735)* ; 1862(899)
g851 and 1859(547)* 1856(417)* 1853(735)* ; 1866(900)
g852 and 1258(674) 432(99) ; 1266(901)
g853 and 1276(595) 432(99) ; 1284(902)
g854 and 1294(612) 432(99) ; 1302(903)
g855 and 1312(693) 432(99) ; 1320(904)
g856 and 1330(710) 432(99) ; 1338(905)
g857 and 1348(631) 432(99) ; 1356(906)
g858 and 1366(648) 432(99) ; 1374(907)
g859 and 980(200) 902(729) ; 983(908)
g860 and 1008(204) 911(724) ; 1011(909)
g861 and 942(441) 649(723) ; 947(910)
g862 and 1510(750)* 1509(752)* 1508(755)* 1507(759)* 1506(764)* 1505(770)* 1504(777)* 1503(749)* ; 1511(911)
g863 and 1493(753)* 1492(756)* 1491(760)* 1490(765)* 1489(771)* 1488(778)* 1487(844)* 1486(751)* ; 1494(912)
g864 and 1476(757)* 1475(761)* 1474(766)* 1473(772)* 1472(779)* 1471(843)* 1470(853)* 1469(754)* ; 1477(913)
g865 and 1459(762)* 1458(767)* 1457(773)* 1456(780)* 1455(842)* 1454(852)* 1453(861)* 1452(758)* ; 1460(914)
g866 and 1442(768)* 1441(774)* 1440(781)* 1439(841)* 1438(851)* 1437(860)* 1436(870)* 1435(763)* ; 1443(915)
g867 and 1425(775)* 1424(782)* 1423(840)* 1422(850)* 1421(859)* 1420(869)* 1419(879)* 1418(769)* ; 1426(916)
g868 and 1408(783)* 1407(839)* 1406(849)* 1405(858)* 1404(868)* 1403(878)* 1402(889)* 1401(776)* ; 1409(917)
g869 and 1391(838)* 1390(848)* 1389(857)* 1388(867)* 1387(877)* 1386(888)* 1385(898)* 1384(784)* ; 1392(918)
g870 and 2237(785) ; 2242(919)
g871 and 2237(785) ; 2245(920)
g872 and 2237(785) ; 2477(921)
g873 and 2185(786) ; 2190(922)
g874 and 2185(786) ; 2193(923)
g875 and 2185(786) ; 2476(924)
g876 and 2132(787) ; 2137(925)
g877 and 2132(787) ; 2140(926)
g878 and 2132(787) ; 2475(927)
g879 and 2080(788) ; 2085(928)
g880 and 2080(788) ; 2088(929)
g881 and 2080(788) ; 2474(930)
g882 and 2025(789) ; 2028(931)
g883 and 2025(789) ; 2031(932)
g884 and 1975(790) ; 1978(933)
g885 and 1975(790) ; 1981(934)
g886 and 1924(791) ; 1927(935)
g887 and 1924(791) ; 1930(936)
g888 and 1874(792) ; 1877(937)
g889 and 1874(792) ; 1880(938)
g890 and 576(793) ; 579(939)
g891 and 360(794) 359(587) ; 361(940)
g892 and 566(797) 565(795) ; 567(941)
g893 and 570(798) 569(796) ; 571(942)
g894 and 2173(845) 2298(237) ; 2383(943)
g895 and 2225(835) 2298(237) ; 2391(944)
g896 and 1963(881) 2289(239) ; 2341(945)
g897 and 2013(871) 2289(239) ; 2354(946)
g898 and 2068(862) 2289(239) ; 2367(947)
g899 and 1862(899) 2285(241) ; 2320(948)
g900 and 2481(150) 2237(785) 2185(786) 2132(787) 2080(788) ; 2482(949)
g901 and 1374(907)* 1373(897)* 1372(887)* 1371(876)* 1370(866)* 1369(856)* 1368(847)* 1367(799)* ; 1375(950)
g902 and 1357(800)* 1356(906)* 1355(896)* 1354(886)* 1353(875)* 1352(865)* 1351(855)* 1350(807)* ; 1358(951)
g903 and 1340(808)* 1339(801)* 1338(905)* 1337(895)* 1336(885)* 1335(874)* 1334(864)* 1333(814)* ; 1341(952)
g904 and 1323(815)* 1322(809)* 1321(802)* 1320(904)* 1319(894)* 1318(884)* 1317(873)* 1316(820)* ; 1324(953)
g905 and 1306(821)* 1305(816)* 1304(810)* 1303(803)* 1302(903)* 1301(893)* 1300(883)* 1299(825)* ; 1307(954)
g906 and 1289(826)* 1288(822)* 1287(817)* 1286(811)* 1285(804)* 1284(902)* 1283(892)* 1282(829)* ; 1290(955)
g907 and 1272(830)* 1271(827)* 1270(823)* 1269(818)* 1268(812)* 1267(805)* 1266(901)* 1265(832)* ; 1273(956)
g908 and 1255(833)* 1254(831)* 1253(828)* 1252(824)* 1251(819)* 1250(813)* 1249(806)* 1248(834)* ; 1256(957)
g909 and 985(378)* 984(408)* 983(908)* ; 986(958)
g910 and 2229(836) ; 2256(959)
g911 and 596(854) 595(837) ; 597(960)
g912 and 2177(846) ; 2204(961)
g913 and 1013(403)* 1012(386)* 1011(909)* ; 1014(962)
g914 and 2072(863) ; 2099(963)
g915 and 2017(872) ; 2042(964)
g916 and 590(891) 589(880) ; 591(965)
g917 and 1967(882) ; 1992(966)
g918 and 1866(900) ; 1891(967)
g919 and 610(432) 576(793) ; 614(968)
g920 and 941(333) 645(890) ; 944(969)
g921 and 579(939) ; 2994(970)
g922 and 579(939) ; 3002(971)
g923 and 567(941) ; 568(972)
g924 and 571(942) ; 2991(973)
g925 and 571(942) ; 2999(974)
g926 and 2383(943) ; 3224(975)
g927 and 2383(943) ; 3232(976)
g928 and 2391(944) ; 3240(977)
g929 and 2391(944) ; 3248(978)
g930 and 2341(945) ; 3158(979)
g931 and 2341(945) ; 3166(980)
g932 and 2354(946) ; 3174(981)
g933 and 2354(946) ; 3182(982)
g934 and 2367(947) ; 3190(983)
g935 and 2367(947) ; 3200(984)
g936 and 2320(948) ; 3124(985)
g937 and 2320(948) ; 3134(986)
g938 and 2242(919) 2229(836) 200(25) ; 2255(987)
g939 and 2190(922) 2177(846) 200(25) ; 2203(988)
g940 and 2085(928) 2072(863) 200(25) ; 2098(989)
g941 and 2028(931) 2017(872) 200(25) ; 2041(990)
g942 and 1978(933) 1967(882) 200(25) ; 1991(991)
g943 and 1877(937) 1866(900) 200(25) ; 1890(992)
g944 and 2245(920) 2229(836) 190(24) ; 2254(993)
g945 and 2193(923) 2177(846) 190(24) ; 2202(994)
g946 and 2088(929) 2072(863) 190(24) ; 2097(995)
g947 and 2031(932) 2017(872) 190(24) ; 2040(996)
g948 and 1981(934) 1967(882) 190(24) ; 1990(997)
g949 and 1880(938) 1866(900) 190(24) ; 1889(998)
g950 and 2478(64) 2477(921) 2476(924) 2475(927) 2474(930) ; 2483(999)
g951 and 2245(920) 2225(835) 179(23) ; 2251(1000)
g952 and 2193(923) 2173(845) 179(23) ; 2199(1001)
g953 and 2088(929) 2068(862) 179(23) ; 2094(1002)
g954 and 2031(932) 2013(871) 179(23) ; 2037(1003)
g955 and 1981(934) 1963(881) 179(23) ; 1987(1004)
g956 and 1880(938) 1862(899) 179(23) ; 1886(1005)
g957 and 2242(919) 2225(835) 169(22) ; 2248(1006)
g958 and 2190(922) 2173(845) 169(22) ; 2196(1007)
g959 and 2085(928) 2068(862) 169(22) ; 2091(1008)
g960 and 2028(931) 2013(871) 169(22) ; 2034(1009)
g961 and 1978(933) 1963(881) 169(22) ; 1984(1010)
g962 and 1877(937) 1862(899) 169(22) ; 1883(1011)
g963 and 597(960) ; 600(1012)
g964 and 591(965) ; 3063(1013)
g965 and 591(965) ; 3071(1014)
g966 and 678(275) 591(965) ; 679(1015)
g967 and 1533(421) 1256(957) ; 1536(1016)
g968 and 617(536)* 616(424)* 614(968)* ; 618(1017)
g969 and 1534(431) 1392(918) ; 1537(1018)
g970 and 665(433) 597(960) ; 669(1019)
g971 and 1581(304) 1273(956) ; 1582(1020)
g972 and 1512(193) 1409(917) ; 1583(1021)
g973 and 1585(305) 1290(955) ; 1586(1022)
g974 and 1512(193) 1426(916) ; 1587(1023)
g975 and 1589(306) 1307(954) ; 1590(1024)
g976 and 1512(193) 1443(915) ; 1591(1025)
g977 and 1593(307) 1324(953) ; 1594(1026)
g978 and 1512(193) 1460(914) ; 1595(1027)
g979 and 1597(308) 1341(952) ; 1598(1028)
g980 and 1512(193) 1477(913) ; 1599(1029)
g981 and 1601(309) 1358(951) ; 1602(1030)
g982 and 1512(193) 1494(912) ; 1603(1031)
g983 and 1605(310) 1375(950) ; 1606(1032)
g984 and 1512(193) 1511(911) ; 1607(1033)
g985 and 1901(336) 986(958) ; 1903(1034)
g986 and 2109(340) 1014(962) ; 2111(1035)
g987 and 2994(970) ; 2998(1036)
g988 and 3002(971) ; 3006(1037)
g989 and 2991(973) ; 2997(1038)
g990 and 2999(974) ; 3005(1039)
g991 and 3224(975) ; 3228(1040)
g992 and 3232(976) ; 3236(1041)
g993 and 3240(977) ; 3244(1042)
g994 and 3248(978) ; 3252(1043)
g995 and 3158(979) ; 3162(1044)
g996 and 3166(980) ; 3170(1045)
g997 and 3174(981) ; 3178(1046)
g998 and 3182(982) ; 3186(1047)
g999 and 3190(983) ; 3194(1048)
g1000 and 3200(984) ; 3204(1049)
g1001 and 3124(985) ; 3128(1050)
g1002 and 3134(986) ; 3138(1051)
g1003 and 2483(999)* 2482(949)* ; 2484(1052)
g1004 and 2251(1000)* 2248(1006)* ; 2257(1053)
g1005 and 2251(1000)* 2248(1006)* ; 2260(1054)
g1006 and 2199(1001)* 2196(1007)* ; 2205(1055)
g1007 and 2199(1001)* 2196(1007)* ; 2208(1056)
g1008 and 2094(1002)* 2091(1008)* ; 2100(1057)
g1009 and 2094(1002)* 2091(1008)* ; 2101(1058)
g1010 and 2037(1003)* 2034(1009)* ; 2043(1059)
g1011 and 2037(1003)* 2034(1009)* ; 2046(1060)
g1012 and 1987(1004)* 1984(1010)* ; 1993(1061)
g1013 and 1987(1004)* 1984(1010)* ; 1996(1062)
g1014 and 1886(1005)* 1883(1011)* ; 1892(1063)
g1015 and 1886(1005)* 1883(1011)* ; 1893(1064)
g1016 and 2256(959)* 2255(987)* 2254(993)* ; 2261(1065)
g1017 and 600(1012) ; 3066(1066)
g1018 and 600(1012) ; 3074(1067)
g1019 and 2204(961)* 2203(988)* 2202(994)* ; 2209(1068)
g1020 and 2117(531)* 2114(388)* 2111(1035)* ; 2120(1069)
g1021 and 2117(531)* 2114(388)* 2111(1035)* ; 2124(1070)
g1022 and 2099(963)* 2098(989)* 2097(995)* ; 2102(1071)
g1023 and 2042(964)* 2041(990)* 2040(996)* ; 2047(1072)
g1024 and 3063(1013) ; 3069(1073)
g1025 and 3071(1014) ; 3077(1074)
g1026 and 1992(966)* 1991(991)* 1990(997)* ; 1997(1075)
g1027 and 1909(545)* 1906(411)* 1903(1034)* ; 1912(1076)
g1028 and 1909(545)* 1906(411)* 1903(1034)* ; 1916(1077)
g1029 and 1891(967)* 1890(992)* 1889(998)* ; 1894(1078)
g1030 and 1538(548)* 1537(1018)* 1536(1016)* ; 1539(1079)
g1031 and 660(274) 568(972) ; 661(1080)
g1032 and 680(420)* 679(1015)* ; 681(1081)
g1033 and 672(533)* 671(426)* 669(1019)* ; 673(1082)
g1034 and 1583(1021)* 1582(1020)* ; 1584(1083)
g1035 and 1587(1023)* 1586(1022)* ; 1588(1084)
g1036 and 1591(1025)* 1590(1024)* ; 1592(1085)
g1037 and 1595(1027)* 1594(1026)* ; 1596(1086)
g1038 and 1599(1029)* 1598(1028)* ; 1600(1087)
g1039 and 1603(1031)* 1602(1030)* ; 1604(1088)
g1040 and 1607(1033)* 1606(1032)* ; 1608(1089)
g1041 and 1647(551) 618(1017) ; 1652(1090)
g1042 and 2997(1038) 2994(970) ; 619(1091)
g1043 and 3005(1039) 3002(971) ; 582(1092)
g1044 and 2998(1036) 2991(973) ; 620(1093)
g1045 and 3006(1037) 2999(974) ; 583(1094)
g1046 and 2302(236) 2205(1055) ; 2455(1095)
g1047 and 2302(236) 2257(1053) ; 2458(1096)
g1048 and 2120(1069) 2298(237) ; 2375(1097)
g1049 and 2293(238) 1993(1061) ; 2445(1098)
g1050 and 2293(238) 2043(1059) ; 2448(1099)
g1051 and 2488(503) 2484(1052) ; 2489(1100)
g1052 and 1912(1076) 2285(241) ; 2328(1101)
g1053 and 2137(925) 2124(1070) 200(25) ; 2150(1102)
g1054 and 1927(935) 1916(1077) 200(25) ; 1940(1103)
g1055 and 2140(926) 2124(1070) 190(24) ; 2149(1104)
g1056 and 1930(936) 1916(1077) 190(24) ; 1939(1105)
g1057 and 2261(1065) 2260(1054) ; 2262(1106)
g1058 and 2209(1068) 2208(1056) ; 2210(1107)
g1059 and 2140(926) 2120(1069) 179(23) ; 2146(1108)
g1060 and 2100(1057) ; 2311(1109)
g1061 and 2102(1071) 2101(1058) ; 2103(1110)
g1062 and 2047(1072) 2046(1060) ; 2048(1111)
g1063 and 1997(1075) 1996(1062) ; 1998(1112)
g1064 and 1930(936) 1912(1076) 179(23) ; 1936(1113)
g1065 and 1892(1063) ; 2271(1114)
g1066 and 1894(1078) 1893(1064) ; 1895(1115)
g1067 and 2137(925) 2120(1069) 169(22) ; 2143(1116)
g1068 and 1927(935) 1912(1076) 169(22) ; 1933(1117)
g1069 and 3069(1073) 3066(1066) ; 606(1118)
g1070 and 3066(1066) ; 3070(1119)
g1071 and 3077(1074) 3074(1067) ; 603(1120)
g1072 and 3074(1067) ; 3078(1121)
g1073 and 2124(1070) ; 2151(1122)
g1074 and 1916(1077) ; 1941(1123)
g1075 and 662(550)* 661(1080)* ; 663(1124)
g1076 and 683(434) 681(1081) ; 689(1125)
g1077 and 1656(552) 673(1082) ; 1661(1126)
g1078 and 1609(577) 1539(1079) ; 1612(1127)
g1079 and 1618(578) 1584(1083) ; 1621(1128)
g1080 and 1627(579) 1588(1084) ; 1630(1129)
g1081 and 1636(580) 1592(1085) ; 1639(1130)
g1082 and 1645(581) 1596(1086) ; 1648(1131)
g1083 and 1654(582) 1600(1087) ; 1657(1132)
g1084 and 1663(583) 1604(1088) ; 1666(1133)
g1085 and 1672(584) 1608(1089) ; 1675(1134)
g1086 and 620(1093) 619(1091) ; 356(1135)
g1087 and 583(1094) 582(1092) ; 357(1136)
g1088 and 2458(1096) ; 2461(1137)
g1089 and 2458(1096) ; 3323(1138)
g1090 and 2375(1097) ; 3208(1139)
g1091 and 2375(1097) ; 3216(1140)
g1092 and 2445(1098) ; 2530(1141)
g1093 and 2448(1099) ; 2451(1142)
g1094 and 2328(1101) ; 3142(1143)
g1095 and 2328(1101) ; 3150(1144)
g1096 and 2151(1122)* 2150(1102)* 2149(1104)* ; 2156(1145)
g1097 and 1941(1123)* 1940(1103)* 1939(1105)* ; 1946(1146)
g1098 and 2262(1106) ; 2388(1147)
g1099 and 2210(1107) ; 2380(1148)
g1100 and 2146(1108)* 2143(1116)* ; 2152(1149)
g1101 and 2146(1108)* 2143(1116)* ; 2155(1150)
g1102 and 2103(1110) ; 2364(1151)
g1103 and 2048(1111) ; 2351(1152)
g1104 and 1998(1112) ; 2338(1153)
g1105 and 1936(1113)* 1933(1117)* ; 1942(1154)
g1106 and 1936(1113)* 1933(1117)* ; 1945(1155)
g1107 and 1895(1115) ; 2317(1156)
g1108 and 691(524)* 690(535)* 689(1125)* ; 692(1157)
g1109 and 3070(1119) 3063(1013) ; 607(1158)
g1110 and 3078(1121) 3071(1014) ; 604(1159)
g1111 and 694(435) 663(1124) ; 700(1160)
g1112 and 357(1136) 356(1135) ; 358(1161)
g1113 and 3323(1138) ; 3329(1162)
g1114 and 3208(1139) ; 3212(1163)
g1115 and 3216(1140) ; 3220(1164)
g1116 and 2293(238) 2152(1149) ; 2454(1165)
g1117 and 2288(240) 1942(1154) ; 2444(1166)
g1118 and 3142(1143) ; 3146(1167)
g1119 and 3150(1144) ; 3154(1168)
g1120 and 2156(1145) 2155(1150) ; 2157(1169)
g1121 and 1946(1146) 1945(1155) ; 1947(1170)
g1122 and 2388(1147) ; 3237(1171)
g1123 and 2388(1147) ; 3245(1172)
g1124 and 2380(1148) ; 3221(1173)
g1125 and 2380(1148) ; 3229(1174)
g1126 and 2152(1149) 2103(1110) ; 2312(1175)
g1127 and 2364(1151) ; 3187(1176)
g1128 and 2364(1151) ; 3197(1177)
g1129 and 2351(1152) ; 3171(1178)
g1130 and 2351(1152) ; 3179(1179)
g1131 and 2338(1153) ; 3155(1180)
g1132 and 2338(1153) ; 3163(1181)
g1133 and 1942(1154) 1895(1115) ; 2272(1182)
g1134 and 2317(1156) ; 3121(1183)
g1135 and 2317(1156) ; 3131(1184)
g1136 and 607(1158) 606(1118) ; 608(1185)
g1137 and 604(1159) 603(1120) ; 605(1186)
g1138 and 702(530)* 701(523)* 700(1160)* ; 703(1187)
g1139 and 1674(554) 692(1157) ; 1679(1188)
g1140 and 3228(1040) 3221(1173) ; 2432(1189)
g1141 and 3236(1041) 3229(1174) ; 2387(1190)
g1142 and 3244(1042) 3237(1171) ; 2395(1191)
g1143 and 3252(1043) 3245(1172) ; 2400(1192)
g1144 and 2454(1165) ; 2533(1193)
g1145 and 3162(1044) 3155(1180) ; 2345(1194)
g1146 and 3170(1045) 3163(1181) ; 2350(1195)
g1147 and 3178(1046) 3171(1178) ; 2358(1196)
g1148 and 3186(1047) 3179(1179) ; 2363(1197)
g1149 and 3194(1048) 3187(1176) ; 3196(1198)
g1150 and 3204(1049) 3197(1177) ; 2371(1199)
g1151 and 2444(1166) ; 2523(1200)
g1152 and 3128(1050) 3121(1183) ; 3130(1201)
g1153 and 3138(1051) 3131(1184) ; 2324(1202)
g1154 and 2157(1169) ; 2372(1203)
g1155 and 1947(1170) ; 2325(1204)
g1156 and 2103(1110) 2210(1107) 2157(1169) 2257(1053) ; 2314(1205)
g1157 and 2262(1106) 2210(1107) 2157(1169) 2103(1110) ; 2309(1206)
g1158 and 3237(1171) ; 3243(1207)
g1159 and 3245(1172) ; 3251(1208)
g1160 and 2205(1055) 2157(1169) 2103(1110) ; 2313(1209)
g1161 and 3221(1173) ; 3227(1210)
g1162 and 3229(1174) ; 3235(1211)
g1163 and 3187(1176) ; 3193(1212)
g1164 and 3197(1177) ; 3203(1213)
g1165 and 1895(1115) 1998(1112) 1947(1170) 2043(1059) ; 2274(1214)
g1166 and 2048(1111) 1998(1112) 1947(1170) 1895(1115) ; 2265(1215)
g1167 and 3171(1178) ; 3177(1216)
g1168 and 3179(1179) ; 3185(1217)
g1169 and 1993(1061) 1947(1170) 1895(1115) ; 2273(1218)
g1170 and 3155(1180) ; 3161(1219)
g1171 and 3163(1181) ; 3169(1220)
g1172 and 3121(1183) ; 3127(1221)
g1173 and 3131(1184) ; 3137(1222)
g1174 and 608(1185) ; 350(1223)
g1175 and 605(1186) ; 349(1224)
g1176 and 1665(553) 703(1187) ; 1670(1225)
g1177 and 3227(1210) 3224(975) ; 2431(1226)
g1178 and 3235(1211) 3232(976) ; 2386(1227)
g1179 and 3243(1207) 3240(977) ; 2394(1228)
g1180 and 3251(1208) 3248(978) ; 2399(1229)
g1181 and 2485(369) 2309(1206) ; 2490(1230)
g1182 and 3161(1219) 3158(979) ; 2344(1231)
g1183 and 3169(1220) 3166(980) ; 2349(1232)
g1184 and 3177(1216) 3174(981) ; 2357(1233)
g1185 and 3185(1217) 3182(982) ; 2362(1234)
g1186 and 3193(1212) 3190(983) ; 3195(1235)
g1187 and 3203(1213) 3200(984) ; 2370(1236)
g1188 and 3127(1221) 3124(985) ; 3129(1237)
g1189 and 3137(1222) 3134(986) ; 2323(1238)
g1190 and 2372(1203) ; 3205(1239)
g1191 and 2372(1203) ; 3213(1240)
g1192 and 2325(1204) ; 3139(1241)
g1193 and 2325(1204) ; 3147(1242)
g1194 and 2265(1215) 2309(1206) ; 372(1243)
g1195 and 2314(1205) 2313(1209) 2312(1175) 2311(1109) ; 2315(1244)
g1196 and 2265(1215) ; 2268(1245)
g1197 and 2274(1214) 2273(1218) 2272(1182) 2271(1114) ; 2275(1246)
g1198 and 350(1223) 349(1224) ; 351(1247)
g1199 and 2302(236) 2315(1244) ; 2464(1248)
g1200 and 3212(1163) 3205(1239) ; 2425(1249)
g1201 and 3220(1164) 3213(1240) ; 2379(1250)
g1202 and 2432(1189) 2431(1226) ; 2433(1251)
g1203 and 2387(1190) 2386(1227) ; 1669(1252)
g1204 and 2395(1191) 2394(1228) ; 2396(1253)
g1205 and 2400(1192) 2399(1229) ; 1678(1254)
g1206 and 2490(1230)* 2489(1100)* ; 2491(1255)
g1207 and 2345(1194) 2344(1231) ; 2346(1256)
g1208 and 2350(1195) 2349(1232) ; 1633(1257)
g1209 and 2358(1196) 2357(1233) ; 2359(1258)
g1210 and 2363(1197) 2362(1234) ; 1642(1259)
g1211 and 3196(1198) 3195(1235) ; 3308(1260)
g1212 and 2371(1199) 2370(1236) ; 1651(1261)
g1213 and 3130(1201) 3129(1237) ; 3272(1262)
g1214 and 2324(1202) 2323(1238) ; 1615(1263)
g1215 and 3146(1167) 3139(1241) ; 2332(1264)
g1216 and 3154(1168) 3147(1242) ; 2337(1265)
g1217 and 3205(1239) ; 3211(1266)
g1218 and 3213(1240) ; 3219(1267)
g1219 and 3139(1241) ; 3145(1268)
g1220 and 3147(1242) ; 3153(1269)
g1221 and 2315(1244) 2265(1215) ; 2307(1270)
g1222 and 2275(1246) ; 2308(1271)
g1223 and 2396(1253) 330(46) ; 2612(1272)
g1224 and 2491(1255) 330(46) ; 3374(1273)
g1225 and 2461(1137) 2433(1251) ; 2518(1274)
g1226 and 2464(1248) ; 2467(1275)
g1227 and 2464(1248) ; 3295(1276)
g1228 and 3211(1266) 3208(1139) ; 2424(1277)
g1229 and 3219(1267) 3216(1140) ; 2378(1278)
g1230 and 2433(1251) ; 3326(1279)
g1231 and 1669(1252) ; 1667(1280)
g1232 and 2396(1253) ; 2439(1281)
g1233 and 1678(1254) ; 1676(1282)
g1234 and 2491(1255) ; 2495(1283)
g1235 and 2346(1256) ; 2406(1284)
g1236 and 2346(1256) ; 2409(1285)
g1237 and 1633(1257) ; 1631(1286)
g1238 and 2359(1258) ; 2415(1287)
g1239 and 2359(1258) ; 2419(1288)
g1240 and 1642(1259) ; 1640(1289)
g1241 and 3308(1260) ; 3312(1290)
g1242 and 1651(1261) ; 1649(1291)
g1243 and 3272(1262) ; 3276(1292)
g1244 and 1615(1263) ; 1613(1293)
g1245 and 3145(1268) 3142(1143) ; 2331(1294)
g1246 and 3153(1269) 3150(1144) ; 2336(1295)
g1247 and 2308(1271) 2307(1270) ; 368(1296)
g1248 and 2612(1272) ; 3406(1297)
g1249 and 2612(1272) ; 3414(1298)
g1250 and 3374(1273) ; 3378(1299)
g1251 and 2518(1274)* 2455(1095)* ; 2519(1300)
g1252 and 3329(1162) 3326(1279) ; 2607(1301)
g1253 and 2415(1287) 2467(1275) ; 2517(1302)
g1254 and 2467(1275) 2419(1288) 2409(1285) ; 2532(1303)
g1255 and 2467(1275) ; 2642(1304)
g1256 and 2467(1275) ; 2645(1305)
g1257 and 3295(1276) ; 3301(1306)
g1258 and 2425(1249) 2424(1277) ; 2426(1307)
g1259 and 2379(1250) 2378(1278) ; 1660(1308)
g1260 and 2433(1251) 2439(1281) ; 2514(1309)
g1261 and 3326(1279) ; 3330(1310)
g1262 and 2439(1281) 2439(1281) ; 3422(1311)
g1263 and 2451(1142) 2409(1285) ; 2531(1312)
g1264 and 2409(1285) 2419(1288) 2495(1283) ; 2511(1313)
g1265 and 2415(1287) 2495(1283) ; 2512(1314)
g1266 and 2409(1285) ; 3290(1315)
g1267 and 2415(1287) ; 3298(1316)
g1268 and 2332(1264) 2331(1294) ; 2333(1317)
g1269 and 2337(1265) 2336(1295) ; 1624(1318)
g1270 and 2268(1245) 2467(1275) ; 2500(1319)
g1271 and 2268(1245) 2495(1283) ; 2505(1320)
g1272 and 368(1296) ; 369(1321)
g1273 and 1646(436) 1649(1291) ; 1650(1322)
g1274 and 1664(438) 1667(1280) ; 1668(1323)
g1275 and 1673(439) 1676(1282) ; 1677(1324)
g1276 and 1610(446) 1613(1293) ; 1614(1325)
g1277 and 1628(448) 1631(1286) ; 1632(1326)
g1278 and 1637(449) 1640(1289) ; 1641(1327)
g1279 and 2642(1304) 2491(1255) 330(46) ; 2643(1328)
g1280 and 3425(130) 3422(1311) ; 2624(1329)
g1281 and 3406(1297) ; 3410(1330)
g1282 and 3414(1298) ; 3418(1331)
g1283 and 2514(1309) 330(46) ; 3398(1332)
g1284 and 2512(1314) 330(46) ; 2567(1333)
g1285 and 2511(1313) 330(46) ; 3350(1334)
g1286 and 2455(1095) 2426(1307) ; 2534(1335)
g1287 and 2519(1300) ; 3313(1336)
g1288 and 2519(1300) ; 2654(1337)
g1289 and 2461(1137) 2433(1251) 2426(1307) ; 2535(1338)
g1290 and 3330(1310) 3323(1138) ; 2608(1339)
g1291 and 3301(1306) 3298(1316) ; 3303(1340)
g1292 and 2426(1307) ; 3316(1341)
g1293 and 1660(1308) ; 1658(1342)
g1294 and 2426(1307) 2433(1251) 2439(1281) ; 2513(1343)
g1295 and 3422(1311) ; 3426(1344)
g1296 and 2532(1303) 2531(1312) 2530(1141) ; 3277(1345)
g1297 and 2517(1302)* 2448(1099)* ; 3287(1346)
g1298 and 3290(1315) ; 3294(1347)
g1299 and 3298(1316) ; 3302(1348)
g1300 and 2333(1317) ; 3280(1349)
g1301 and 2333(1317) ; 2401(1350)
g1302 and 1624(1318) ; 1622(1351)
g1303 and 2505(1320) ; 3253(1352)
g1304 and 2500(1319)* 2275(1246)* ; 2501(1353)
g1305 and 1643(727)* 1641(1327)* 1639(1130)* ; 1644(1354)
g1306 and 1634(730)* 1632(1326)* 1630(1129)* ; 1635(1355)
g1307 and 1616(733)* 1614(1325)* 1612(1127)* ; 1617(1356)
g1308 and 1652(1090)* 1650(1322)* 1648(1131)* ; 1653(1357)
g1309 and 1670(1225)* 1668(1323)* 1666(1133)* ; 1671(1358)
g1310 and 1679(1188)* 1677(1324)* 1675(1134)* ; 1680(1359)
g1311 and 3426(1344) 3419(51) ; 2625(1360)
g1312 and 3398(1332) ; 3402(1361)
g1313 and 2513(1343) 330(46) ; 2589(1362)
g1314 and 2567(1333) ; 3358(1363)
g1315 and 2567(1333) ; 3366(1364)
g1316 and 3350(1334) ; 3354(1365)
g1317 and 2654(1337) 2519(1300) ; 398(1366)
g1318 and 3313(1336) ; 3319(1367)
g1319 and 2654(1337) ; 2657(1368)
g1320 and 2608(1339) 2607(1301) ; 2609(1369)
g1321 and 2467(1275) 2419(1288) 2406(1284) 2401(1350) ; 2526(1370)
g1322 and 2645(1305)* 2643(1328)* ; 932(1371)
g1323 and 2645(1305)* 2643(1328)* ; 2647(1372)
g1324 and 3302(1348) 3295(1276) ; 3304(1373)
g1325 and 3316(1341) ; 3320(1374)
g1326 and 2445(1098) 2401(1350) ; 2524(1375)
g1327 and 3277(1345) ; 3283(1376)
g1328 and 2451(1142) 2406(1284) 2401(1350) ; 2525(1377)
g1329 and 3294(1347) 3287(1346) ; 2563(1378)
g1330 and 3287(1346) ; 3293(1379)
g1331 and 2535(1338) 2534(1335) 2533(1193) ; 3305(1380)
g1332 and 2419(1288) 2409(1285) 2401(1350) 2495(1283) ; 2508(1381)
g1333 and 3280(1349) ; 3284(1382)
g1334 and 3253(1352) ; 3259(1383)
g1335 and 2501(1353) ; 3264(1384)
g1336 and 2501(1353) ; 2629(1385)
g1337 and 1655(437) 1658(1342) ; 1659(1386)
g1338 and 1619(447) 1622(1351) ; 1623(1387)
g1339 and 2680(568) 1617(1356) ; 2687(1388)
g1340 and 2718(570) 1635(1355) ; 2725(1389)
g1341 and 2735(571) 1644(1354) ; 2742(1390)
g1342 and 2753(572) 1653(1357) ; 2760(1391)
g1343 and 2787(574) 1671(1358) ; 2794(1392)
g1344 and 2804(575) 1680(1359) ; 2811(1393)
g1345 and 2657(1368) 2514(1309) 330(46) ; 397(1394)
g1346 and 2625(1360) 2624(1329) ; 2626(1395)
g1347 and 2589(1362) ; 3382(1396)
g1348 and 2589(1362) ; 3390(1397)
g1349 and 3358(1363) ; 3362(1398)
g1350 and 3366(1364) ; 3370(1399)
g1351 and 2508(1381) 330(46) ; 2544(1400)
g1352 and 3320(1374) 3313(1336) ; 3322(1401)
g1353 and 2609(1369) ; 3403(1402)
g1354 and 2609(1369) ; 3411(1403)
g1355 and 2647(1372) ; 2650(1404)
g1356 and 3304(1373) 3303(1340) ; 3371(1405)
g1357 and 3319(1367) 3316(1341) ; 3321(1406)
g1358 and 3284(1382) 3277(1345) ; 3286(1407)
g1359 and 3305(1380) ; 3311(1408)
g1360 and 2508(1381) ; 3256(1409)
g1361 and 3293(1379) 3290(1315) ; 2562(1410)
g1362 and 3312(1290) 3305(1380) ; 2585(1411)
g1363 and 2526(1370) 2525(1377) 2524(1375) 2523(1200) ; 2527(1412)
g1364 and 3283(1376) 3280(1349) ; 3285(1413)
g1365 and 3264(1384) ; 3268(1414)
g1366 and 2629(1385) ; 2632(1415)
g1367 and 2629(1385) 2501(1353) ; 2634(1416)
g1368 and 1625(732)* 1623(1387)* 1621(1128)* ; 1626(1417)
g1369 and 1661(1126)* 1659(1386)* 1657(1132)* ; 1662(1418)
g1370 and 927(347) 932(1371) ; 933(1419)
g1371 and 2632(1415) 2505(1320) 330(46) ; 2633(1420)
g1372 and 3410(1330) 3403(1402) ; 2616(1421)
g1373 and 3418(1331) 3411(1403) ; 2622(1422)
g1374 and 3382(1396) ; 3386(1423)
g1375 and 3390(1397) ; 3394(1424)
g1376 and 3378(1299) 3371(1405) ; 2580(1425)
g1377 and 2544(1400) ; 3334(1426)
g1378 and 2544(1400) ; 3342(1427)
g1379 and 398(1366)* 397(1394)* ; 399(1428)
g1380 and 3322(1401) 3321(1406) ; 3395(1429)
g1381 and 3403(1402) ; 3409(1430)
g1382 and 3411(1403) ; 3417(1431)
g1383 and 2650(1404) ; 3454(1432)
g1384 and 3371(1405) ; 3377(1433)
g1385 and 3286(1407) 3285(1413) ; 3347(1434)
g1386 and 2563(1378) 2562(1410) ; 2564(1435)
g1387 and 3256(1409) ; 3260(1436)
g1388 and 3311(1408) 3308(1260) ; 2584(1437)
g1389 and 2527(1412) ; 3261(1438)
g1390 and 2527(1412) ; 3269(1439)
g1391 and 3259(1383) 3256(1409) ; 2536(1440)
g1392 and 938(722)* 933(1419)* 929(734)* ; 362(1441)
g1393 and 938(722)* 933(1419)* 929(734)* ; 1030(1442)
g1394 and 2803(562) 2626(1395) ; 2808(1443)
g1395 and 2699(569) 1626(1417) ; 2706(1444)
g1396 and 2770(573) 1662(1418) ; 2777(1445)
g1397 and 2802(469) 2626(1395) ; 2805(1446)
g1398 and 3409(1430) 3406(1297) ; 2615(1447)
g1399 and 3417(1431) 3414(1298) ; 2621(1448)
g1400 and 3402(1361) 3395(1429) ; 2602(1449)
g1401 and 3377(1433) 3374(1273) ; 2579(1450)
g1402 and 3354(1365) 3347(1434) ; 2557(1451)
g1403 and 3334(1426) ; 3338(1452)
g1404 and 3342(1427) ; 3346(1453)
g1405 and 3395(1429) ; 3401(1454)
g1406 and 3454(1432) ; 3458(1455)
g1407 and 3347(1434) ; 3353(1456)
g1408 and 2564(1435) ; 3355(1457)
g1409 and 2564(1435) ; 3363(1458)
g1410 and 2585(1411) 2584(1437) ; 2586(1459)
g1411 and 3261(1438) ; 3267(1460)
g1412 and 3269(1439) ; 3275(1461)
g1413 and 3276(1292) 3269(1439) ; 2540(1462)
g1414 and 3260(1436) 3253(1352) ; 2537(1463)
g1415 and 3268(1414) 3261(1438) ; 3112(1464)
g1416 and 2634(1416)* 2633(1420)* ; 2635(1465)
g1417 and 1030(1442) ; 363(1466)
g1418 and 2811(1393)* 2808(1443)* 2805(1446)* ; 2814(1467)
g1419 and 2811(1393)* 2808(1443)* 2805(1446)* ; 2816(1468)
g1420 and 2616(1421) 2615(1447) ; 2617(1469)
g1421 and 2622(1422) 2621(1448) ; 2623(1470)
g1422 and 3401(1454) 3398(1332) ; 2601(1471)
g1423 and 2580(1425) 2579(1450) ; 2581(1472)
g1424 and 3362(1398) 3355(1457) ; 2571(1473)
g1425 and 3370(1399) 3363(1458) ; 2577(1474)
g1426 and 3353(1456) 3350(1334) ; 2556(1475)
g1427 and 3355(1457) ; 3361(1476)
g1428 and 3363(1458) ; 3369(1477)
g1429 and 2586(1459) ; 3379(1478)
g1430 and 2586(1459) ; 3387(1479)
g1431 and 3275(1461) 3272(1262) ; 2539(1480)
g1432 and 2537(1463) 2536(1440) ; 2538(1481)
g1433 and 3267(1460) 3264(1384) ; 3111(1482)
g1434 and 2635(1465) ; 2638(1483)
g1435 and 363(1466) 362(1441) ; 364(1484)
g1436 and 2814(1467) ; 3459(1485)
g1437 and 2816(1468) ; 395(1486)
g1438 and 2623(1470) ; 3451(1487)
g1439 and 2602(1449) 2601(1471) ; 2603(1488)
g1440 and 3386(1423) 3379(1478) ; 2593(1489)
g1441 and 3394(1424) 3387(1479) ; 2598(1490)
g1442 and 3361(1476) 3358(1363) ; 2570(1491)
g1443 and 3369(1477) 3366(1364) ; 2576(1492)
g1444 and 2557(1451) 2556(1475) ; 2558(1493)
g1445 and 2538(1481) 330(46) ; 3116(1494)
g1446 and 2647(1372) 2617(1469) ; 3446(1495)
g1447 and 3379(1478) ; 3385(1496)
g1448 and 3387(1479) ; 3393(1497)
g1449 and 2540(1462) 2539(1480) ; 2541(1498)
g1450 and 3112(1464) 3111(1482) ; 3113(1499)
g1451 and 2638(1483) ; 3438(1500)
g1452 and 2734(558) 2581(1472) ; 2739(1501)
g1453 and 2733(465) 2581(1472) ; 2736(1502)
g1454 and 2785(468) 2617(1469) ; 2788(1503)
g1455 and 395(1486) 2814(1467) ; 396(1504)
g1456 and 3459(1485) ; 3465(1505)
g1457 and 3451(1487) ; 3457(1506)
g1458 and 2603(1488) ; 3443(1507)
g1459 and 3385(1496) 3382(1396) ; 2592(1508)
g1460 and 3393(1497) 3390(1397) ; 2597(1509)
g1461 and 2571(1473) 2570(1491) ; 2572(1510)
g1462 and 2577(1474) 2576(1492) ; 2578(1511)
g1463 and 2558(1493) ; 3427(1512)
g1464 and 3116(1494) ; 3120(1513)
g1465 and 3458(1455) 3451(1487) ; 2677(1514)
g1466 and 3446(1495) ; 3450(1515)
g1467 and 2541(1498) ; 3331(1516)
g1468 and 2541(1498) ; 3339(1517)
g1469 and 3113(1499) ; 3119(1518)
g1470 and 3438(1500) ; 3442(1519)
g1471 and 2697(463) 2558(1493) ; 2700(1520)
g1472 and 2742(1390)* 2739(1501)* 2736(1502)* ; 2745(1521)
g1473 and 2742(1390)* 2739(1501)* 2736(1502)* ; 2748(1522)
g1474 and 2768(467) 2603(1488) ; 2771(1523)
g1475 and 3450(1515) 3443(1507) ; 2672(1524)
g1476 and 3443(1507) ; 3449(1525)
g1477 and 2593(1489) 2592(1508) ; 2594(1526)
g1478 and 2598(1490) 2597(1509) ; 2599(1527)
g1479 and 2578(1511) ; 3435(1528)
g1480 and 3427(1512) ; 3433(1529)
g1481 and 3338(1452) 3331(1516) ; 2548(1530)
g1482 and 3346(1453) 3339(1517) ; 2553(1531)
g1483 and 3119(1518) 3116(1494) ; 954(1532)
g1484 and 3457(1506) 3454(1432) ; 2676(1533)
g1485 and 3331(1516) ; 3337(1534)
g1486 and 3339(1517) ; 3345(1535)
g1487 and 3120(1513) 3113(1499) ; 955(1536)
g1488 and 2635(1465) 2572(1510) ; 3430(1537)
g1489 and 2716(464) 2572(1510) ; 2719(1538)
g1490 and 2745(1521) ; 3491(1539)
g1491 and 2745(1521) ; 3499(1540)
g1492 and 2748(1522) ; 383(1541)
g1493 and 2599(1527) ; 2600(1542)
g1494 and 3435(1528) ; 3441(1543)
g1495 and 3433(1529) 3430(1537) ; 2664(1544)
g1496 and 3337(1534) 3334(1426) ; 2547(1545)
g1497 and 3345(1535) 3342(1427) ; 2552(1546)
g1498 and 955(1536) 954(1532) ; 950(1547)
g1499 and 2650(1404) 2594(1526) 2603(1488) 2617(1469) ; 2662(1548)
g1500 and 2677(1514) 2676(1533) ; 2674(1549)
g1501 and 3449(1525) 3446(1495) ; 2671(1550)
g1502 and 3442(1519) 3435(1528) ; 2670(1551)
g1503 and 3430(1537) ; 3434(1552)
g1504 and 383(1541) 2745(1521) ; 384(1553)
g1505 and 3491(1539) ; 3497(1554)
g1506 and 3499(1540) ; 3505(1555)
g1507 and 2751(466) 2594(1526) ; 2754(1556)
g1508 and 2672(1524) 2671(1550) ; 2673(1557)
g1509 and 3434(1552) 3427(1512) ; 2665(1558)
g1510 and 2548(1530) 2547(1545) ; 2549(1559)
g1511 and 2553(1531) 2552(1546) ; 2554(1560)
g1512 and 2650(1404)* 2600(1542)* ; 2661(1561)
g1513 and 2674(1549) ; 2675(1562)
g1514 and 3441(1543) 3438(1500) ; 2669(1563)
g1515 and 943(445) 950(1547) ; 951(1564)
g1516 and 2665(1558) 2664(1544) ; 2666(1565)
g1517 and 2554(1560) ; 2555(1566)
g1518 and 2662(1548)* 2661(1561)* ; 2663(1567)
g1519 and 2638(1483) 2549(1559) 2558(1493) 2572(1510) ; 2659(1568)
g1520 and 2670(1551) 2669(1563) ; 2667(1569)
g1521 and 951(1564)* 947(910)* 944(969)* ; 365(1570)
g1522 and 951(1564)* 947(910)* 944(969)* ; 1031(1571)
g1523 and 2769(560) 2673(1557) ; 2774(1572)
g1524 and 2786(561) 2675(1562) ; 2791(1573)
g1525 and 2678(462) 2549(1559) ; 2681(1574)
g1526 and 2638(1483)* 2555(1566)* ; 2658(1575)
g1527 and 2667(1569) ; 2668(1576)
g1528 and 1031(1571) ; 366(1577)
g1529 and 2698(556) 2666(1565) ; 2703(1578)
g1530 and 2752(559) 2663(1567) ; 2757(1579)
g1531 and 2777(1445)* 2774(1572)* 2771(1523)* ; 2780(1580)
g1532 and 2777(1445)* 2774(1572)* 2771(1523)* ; 2782(1581)
g1533 and 2794(1392)* 2791(1573)* 2788(1503)* ; 2797(1582)
g1534 and 2794(1392)* 2791(1573)* 2788(1503)* ; 2799(1583)
g1535 and 2659(1568)* 2658(1575)* ; 2660(1584)
g1536 and 366(1577) 365(1570) ; 367(1585)
g1537 and 2717(557) 2668(1576) ; 2722(1586)
g1538 and 2706(1444)* 2703(1578)* 2700(1520)* ; 2709(1587)
g1539 and 2706(1444)* 2703(1578)* 2700(1520)* ; 2713(1588)
g1540 and 2760(1391)* 2757(1579)* 2754(1556)* ; 2763(1589)
g1541 and 2760(1391)* 2757(1579)* 2754(1556)* ; 2765(1590)
g1542 and 2780(1580) ; 3467(1591)
g1543 and 2782(1581) ; 389(1592)
g1544 and 2797(1582) ; 3462(1593)
g1545 and 2799(1583) ; 392(1594)
g1546 and 2871(128) 2709(1587) ; 2883(1595)
g1547 and 2679(555) 2660(1584) ; 2684(1596)
g1548 and 2709(1587) 2709(1587) ; 378(1597)
g1549 and 2709(1587) ; 3507(1598)
g1550 and 2725(1389)* 2722(1586)* 2719(1538)* ; 2728(1599)
g1551 and 2725(1389)* 2722(1586)* 2719(1538)* ; 2730(1600)
g1552 and 2763(1589) ; 3470(1601)
g1553 and 2765(1590) ; 386(1602)
g1554 and 389(1592) 2780(1580) ; 390(1603)
g1555 and 3467(1591) ; 3473(1604)
g1556 and 392(1594) 2797(1582) ; 393(1605)
g1557 and 3462(1593) ; 3466(1606)
g1558 and 3465(1505) 3462(1593) ; 2821(1607)
g1559 and 2765(1590) 2782(1581) 2799(1583) 2816(1468) ; 2922(1608)
g1560 and 2883(1595) ; 3544(1609)
g1561 and 2883(1595) ; 3552(1610)
g1562 and 2687(1388)* 2684(1596)* 2681(1574)* ; 2690(1611)
g1563 and 2687(1388)* 2684(1596)* 2681(1574)* ; 2694(1612)
g1564 and 3507(1598) ; 3513(1613)
g1565 and 2728(1599) ; 2839(1614)
g1566 and 2730(1600) ; 380(1615)
g1567 and 386(1602) 2763(1589) ; 387(1616)
g1568 and 3473(1604) 3470(1601) ; 2826(1617)
g1569 and 3470(1601) ; 3474(1618)
g1570 and 3466(1606) 3459(1485) ; 2822(1619)
g1571 and 2690(1611) 2871(128) ; 2880(1620)
g1572 and 3544(1609) ; 3548(1621)
g1573 and 3552(1610) ; 3556(1622)
g1574 and 2874(129) 2694(1612) 2713(1588) ; 2928(1623)
g1575 and 2690(1611) 2690(1611) ; 375(1624)
g1576 and 2690(1611) ; 3510(1625)
g1577 and 380(1615) 2728(1599) ; 381(1626)
g1578 and 2839(1614) ; 3494(1627)
g1579 and 2839(1614) ; 3502(1628)
g1580 and 2694(1612) 2713(1588) 2730(1600) 2748(1522) ; 2925(1629)
g1581 and 3474(1618) 3467(1591) ; 2827(1630)
g1582 and 2822(1619) 2821(1607) ; 2823(1631)
g1583 and 2880(1620) ; 3541(1632)
g1584 and 2880(1620) ; 3549(1633)
g1585 and 3510(1625) ; 3514(1634)
g1586 and 3513(1613) 3510(1625) ; 3515(1635)
g1587 and 3494(1627) ; 3498(1636)
g1588 and 3502(1628) ; 3506(1637)
g1589 and 3497(1554) 3494(1627) ; 2842(1638)
g1590 and 3505(1555) 3502(1628) ; 2852(1639)
g1591 and 2827(1630) 2826(1617) ; 2828(1640)
g1592 and 2823(1631) ; 3475(1641)
g1593 and 2823(1631) ; 3483(1642)
g1594 and 2925(1629) 2922(1608) ; 406(1643)
g1595 and 2925(1629) 2922(1608) ; 2929(1644)
g1596 and 3541(1632) ; 3547(1645)
g1597 and 3549(1633) ; 3555(1646)
g1598 and 3548(1621) 3541(1632) ; 2887(1647)
g1599 and 3556(1622) 3549(1633) ; 2896(1648)
g1600 and 2929(1644)* 2928(1623)* ; 2930(1649)
g1601 and 3514(1634) 3507(1598) ; 3516(1650)
g1602 and 3498(1636) 3491(1539) ; 2843(1651)
g1603 and 3506(1637) 3499(1540) ; 2853(1652)
g1604 and 2828(1640) ; 3478(1653)
g1605 and 2828(1640) ; 3486(1654)
g1606 and 3475(1641) ; 3481(1655)
g1607 and 3483(1642) ; 3489(1656)
g1608 and 406(1643) ; 407(1657)
g1609 and 3547(1645) 3544(1609) ; 2886(1658)
g1610 and 3555(1646) 3552(1610) ; 2895(1659)
g1611 and 2930(1649) 213(26) ; 408(1660)
g1612 and 3516(1650) 3515(1635) ; 3520(1661)
g1613 and 2843(1651) 2842(1638) ; 2844(1662)
g1614 and 2853(1652) 2852(1639) ; 2848(1663)
g1615 and 3481(1655) 3478(1653) ; 2831(1664)
g1616 and 3478(1653) ; 3482(1665)
g1617 and 3489(1656) 3486(1654) ; 2836(1666)
g1618 and 3486(1654) ; 3490(1667)
g1619 and 2887(1647) 2886(1658) ; 2888(1668)
g1620 and 2896(1648) 2895(1659) ; 2891(1669)
g1621 and 408(1660) ; 409(1670)
g1622 and 3520(1661) ; 3524(1671)
g1623 and 2844(1662) ; 3517(1672)
g1624 and 2848(1663) ; 2849(1673)
g1625 and 3482(1665) 3475(1641) ; 2832(1674)
g1626 and 3490(1667) 3483(1642) ; 2837(1675)
g1627 and 2903(349) 2888(1668) 2849(1673) ; 2908(1676)
g1628 and 2900(350) 2888(1668) 2844(1662) ; 2906(1677)
g1629 and 2891(1669) ; 2892(1678)
g1630 and 3524(1671) 3517(1672) ; 2855(1679)
g1631 and 3517(1672) ; 3523(1680)
g1632 and 2832(1674) 2831(1664) ; 2833(1681)
g1633 and 2837(1675) 2836(1666) ; 2838(1682)
g1634 and 2903(349) 2892(1678) 2844(1662) ; 2907(1683)
g1635 and 2900(350) 2892(1678) 2849(1673) ; 2909(1684)
g1636 and 3523(1680) 3520(1661) ; 2854(1685)
g1637 and 2833(1681) ; 3525(1686)
g1638 and 2833(1681) ; 3533(1687)
g1639 and 2838(1682) ; 2913(1688)
g1640 and 2909(1684)* 2908(1676)* 2907(1683)* 2906(1677)* ; 2910(1689)
g1641 and 2855(1679) 2854(1685) ; 2856(1690)
g1642 and 3525(1686) ; 3531(1691)
g1643 and 3533(1687) ; 3539(1692)
g1644 and 2913(1688) ; 3560(1693)
g1645 and 2913(1688) ; 3568(1694)
g1646 and 2910(1689) ; 3557(1695)
g1647 and 2910(1689) ; 3565(1696)
g1648 and 2856(1690) ; 3528(1697)
g1649 and 2856(1690) ; 3536(1698)
g1650 and 3560(1693) ; 3564(1699)
g1651 and 3568(1694) ; 3572(1700)
g1652 and 3564(1699) 3557(1695) ; 2921(1701)
g1653 and 3557(1695) ; 3563(1702)
g1654 and 3572(1700) 3565(1696) ; 2917(1703)
g1655 and 3565(1696) ; 3571(1704)
g1656 and 3528(1697) ; 3532(1705)
g1657 and 3536(1698) ; 3540(1706)
g1658 and 3531(1691) 3528(1697) ; 2863(1707)
g1659 and 3539(1692) 3536(1698) ; 2859(1708)
g1660 and 3532(1705) 3525(1686) ; 2864(1709)
g1661 and 3540(1706) 3533(1687) ; 2860(1710)
g1662 and 3563(1702) 3560(1693) ; 2920(1711)
g1663 and 3571(1704) 3568(1694) ; 2916(1712)
g1664 and 2921(1701) 2920(1711) ; 403(1713)
g1665 and 2917(1703) 2916(1712) ; 404(1714)
g1666 and 2864(1709) 2863(1707) ; 400(1715)
g1667 and 2860(1710) 2859(1708) ; 401(1716)
g1668 and 404(1714) 403(1713) ; 405(1717)
g1669 and 401(1716) 400(1715) ; 402(1718)
g1670 not 257(34) ; 257(34)*
g1671 not 264(35) ; 264(35)*
g1672 not 41(4) ; 41(4)*
g1673 not 45(5) ; 45(5)*
g1674 not 1698(48) ; 1698(48)*
g1675 not 33(3) ; 33(3)*
g1676 not 2865(61) ; 2865(61)*
g1677 not 2868(50) ; 2868(50)*
g1678 not 1032(115) ; 1032(115)*
g1679 not 1035(63) ; 1035(63)*
g1680 not 1540(111) ; 1540(111)*
g1681 not 169(22) ; 169(22)*
g1682 not 758(108) ; 758(108)*
g1683 not 20(2) ; 20(2)*
g1684 not 2051(104) ; 2051(104)*
g1685 not 1(0) ; 1(0)*
g1686 not 1828(110) ; 1828(110)*
g1687 not 1772(212) ; 1772(212)*
g1688 not 116(13) ; 116(13)*
g1689 not 1773(345) ; 1773(345)*
g1690 not 107(12) ; 107(12)*
g1691 not 97(11) ; 97(11)*
g1692 not 87(10) ; 87(10)*
g1693 not 77(9) ; 77(9)*
g1694 not 68(8) ; 68(8)*
g1695 not 58(7) ; 58(7)*
g1696 not 50(6) ; 50(6)*
g1697 not 1768(351) ; 1768(351)*
g1698 not 1769(221) ; 1769(221)*
g1699 not 1770(357) ; 1770(357)*
g1700 not 1761(352) ; 1761(352)*
g1701 not 1762(223) ; 1762(223)*
g1702 not 1763(358) ; 1763(358)*
g1703 not 1754(353) ; 1754(353)*
g1704 not 1755(225) ; 1755(225)*
g1705 not 1756(360) ; 1756(360)*
g1706 not 1747(381) ; 1747(381)*
g1707 not 1748(228) ; 1748(228)*
g1708 not 1749(362) ; 1749(362)*
g1709 not 1740(385) ; 1740(385)*
g1710 not 1741(230) ; 1741(230)*
g1711 not 1742(364) ; 1742(364)*
g1712 not 1733(389) ; 1733(389)*
g1713 not 1734(232) ; 1734(232)*
g1714 not 1735(365) ; 1735(365)*
g1715 not 1726(396) ; 1726(396)*
g1716 not 1727(234) ; 1727(234)*
g1717 not 1728(367) ; 1728(367)*
g1718 not 1719(402) ; 1719(402)*
g1719 not 1720(235) ; 1720(235)*
g1720 not 1721(368) ; 1721(368)*
g1721 not 1025(244) ; 1025(244)*
g1722 not 1026(354) ; 1026(354)*
g1723 not 1027(393) ; 1027(393)*
g1724 not 1004(252) ; 1004(252)*
g1725 not 1005(392) ; 1005(392)*
g1726 not 1006(409) ; 1006(409)*
g1727 not 1018(253) ; 1018(253)*
g1728 not 1019(382) ; 1019(382)*
g1729 not 1020(398) ; 1020(398)*
g1730 not 997(259) ; 997(259)*
g1731 not 998(397) ; 998(397)*
g1732 not 999(415) ; 999(415)*
g1733 not 976(266) ; 976(266)*
g1734 not 977(414) ; 977(414)*
g1735 not 978(379) ; 978(379)*
g1736 not 990(267) ; 990(267)*
g1737 not 991(404) ; 991(404)*
g1738 not 992(418) ; 992(418)*
g1739 not 917(549) ; 917(549)*
g1740 not 920(361) ; 920(361)*
g1741 not 923(482) ; 923(482)*
g1742 not 2234(480) ; 2234(480)*
g1743 not 2235(472) ; 2235(472)*
g1744 not 2236(748) ; 2236(748)*
g1745 not 2182(483) ; 2182(483)*
g1746 not 2183(473) ; 2183(473)*
g1747 not 2184(747) ; 2184(747)*
g1748 not 2129(484) ; 2129(484)*
g1749 not 2130(474) ; 2130(474)*
g1750 not 2131(746) ; 2131(746)*
g1751 not 2077(487) ; 2077(487)*
g1752 not 2078(475) ; 2078(475)*
g1753 not 2079(745) ; 2079(745)*
g1754 not 2022(489) ; 2022(489)*
g1755 not 2023(476) ; 2023(476)*
g1756 not 2024(744) ; 2024(744)*
g1757 not 1972(493) ; 1972(493)*
g1758 not 1973(477) ; 1973(477)*
g1759 not 1974(743) ; 1974(743)*
g1760 not 1921(495) ; 1921(495)*
g1761 not 1922(478) ; 1922(478)*
g1762 not 1923(742) ; 1923(742)*
g1763 not 1871(499) ; 1871(499)*
g1764 not 1872(479) ; 1872(479)*
g1765 not 1873(741) ; 1873(741)*
g1766 not 2216(740) ; 2216(740)*
g1767 not 2219(380) ; 2219(380)*
g1768 not 2222(520) ; 2222(520)*
g1769 not 2164(739) ; 2164(739)*
g1770 not 2167(384) ; 2167(384)*
g1771 not 2170(525) ; 2170(525)*
g1772 not 2059(738) ; 2059(738)*
g1773 not 2062(395) ; 2062(395)*
g1774 not 2065(534) ; 2065(534)*
g1775 not 2004(737) ; 2004(737)*
g1776 not 2007(401) ; 2007(401)*
g1777 not 2010(537) ; 2010(537)*
g1778 not 1954(736) ; 1954(736)*
g1779 not 1957(407) ; 1957(407)*
g1780 not 1960(540) ; 1960(540)*
g1781 not 641(728) ; 641(728)*
g1782 not 644(269) ; 644(269)*
g1783 not 1853(735) ; 1853(735)*
g1784 not 1856(417) ; 1856(417)*
g1785 not 1859(547) ; 1859(547)*
g1786 not 1503(749) ; 1503(749)*
g1787 not 1504(777) ; 1504(777)*
g1788 not 1505(770) ; 1505(770)*
g1789 not 1506(764) ; 1506(764)*
g1790 not 1507(759) ; 1507(759)*
g1791 not 1508(755) ; 1508(755)*
g1792 not 1509(752) ; 1509(752)*
g1793 not 1510(750) ; 1510(750)*
g1794 not 1486(751) ; 1486(751)*
g1795 not 1487(844) ; 1487(844)*
g1796 not 1488(778) ; 1488(778)*
g1797 not 1489(771) ; 1489(771)*
g1798 not 1490(765) ; 1490(765)*
g1799 not 1491(760) ; 1491(760)*
g1800 not 1492(756) ; 1492(756)*
g1801 not 1493(753) ; 1493(753)*
g1802 not 1469(754) ; 1469(754)*
g1803 not 1470(853) ; 1470(853)*
g1804 not 1471(843) ; 1471(843)*
g1805 not 1472(779) ; 1472(779)*
g1806 not 1473(772) ; 1473(772)*
g1807 not 1474(766) ; 1474(766)*
g1808 not 1475(761) ; 1475(761)*
g1809 not 1476(757) ; 1476(757)*
g1810 not 1452(758) ; 1452(758)*
g1811 not 1453(861) ; 1453(861)*
g1812 not 1454(852) ; 1454(852)*
g1813 not 1455(842) ; 1455(842)*
g1814 not 1456(780) ; 1456(780)*
g1815 not 1457(773) ; 1457(773)*
g1816 not 1458(767) ; 1458(767)*
g1817 not 1459(762) ; 1459(762)*
g1818 not 1435(763) ; 1435(763)*
g1819 not 1436(870) ; 1436(870)*
g1820 not 1437(860) ; 1437(860)*
g1821 not 1438(851) ; 1438(851)*
g1822 not 1439(841) ; 1439(841)*
g1823 not 1440(781) ; 1440(781)*
g1824 not 1441(774) ; 1441(774)*
g1825 not 1442(768) ; 1442(768)*
g1826 not 1418(769) ; 1418(769)*
g1827 not 1419(879) ; 1419(879)*
g1828 not 1420(869) ; 1420(869)*
g1829 not 1421(859) ; 1421(859)*
g1830 not 1422(850) ; 1422(850)*
g1831 not 1423(840) ; 1423(840)*
g1832 not 1424(782) ; 1424(782)*
g1833 not 1425(775) ; 1425(775)*
g1834 not 1401(776) ; 1401(776)*
g1835 not 1402(889) ; 1402(889)*
g1836 not 1403(878) ; 1403(878)*
g1837 not 1404(868) ; 1404(868)*
g1838 not 1405(858) ; 1405(858)*
g1839 not 1406(849) ; 1406(849)*
g1840 not 1407(839) ; 1407(839)*
g1841 not 1408(783) ; 1408(783)*
g1842 not 1384(784) ; 1384(784)*
g1843 not 1385(898) ; 1385(898)*
g1844 not 1386(888) ; 1386(888)*
g1845 not 1387(877) ; 1387(877)*
g1846 not 1388(867) ; 1388(867)*
g1847 not 1389(857) ; 1389(857)*
g1848 not 1390(848) ; 1390(848)*
g1849 not 1391(838) ; 1391(838)*
g1850 not 1367(799) ; 1367(799)*
g1851 not 1368(847) ; 1368(847)*
g1852 not 1369(856) ; 1369(856)*
g1853 not 1370(866) ; 1370(866)*
g1854 not 1371(876) ; 1371(876)*
g1855 not 1372(887) ; 1372(887)*
g1856 not 1373(897) ; 1373(897)*
g1857 not 1374(907) ; 1374(907)*
g1858 not 1350(807) ; 1350(807)*
g1859 not 1351(855) ; 1351(855)*
g1860 not 1352(865) ; 1352(865)*
g1861 not 1353(875) ; 1353(875)*
g1862 not 1354(886) ; 1354(886)*
g1863 not 1355(896) ; 1355(896)*
g1864 not 1356(906) ; 1356(906)*
g1865 not 1357(800) ; 1357(800)*
g1866 not 1333(814) ; 1333(814)*
g1867 not 1334(864) ; 1334(864)*
g1868 not 1335(874) ; 1335(874)*
g1869 not 1336(885) ; 1336(885)*
g1870 not 1337(895) ; 1337(895)*
g1871 not 1338(905) ; 1338(905)*
g1872 not 1339(801) ; 1339(801)*
g1873 not 1340(808) ; 1340(808)*
g1874 not 1316(820) ; 1316(820)*
g1875 not 1317(873) ; 1317(873)*
g1876 not 1318(884) ; 1318(884)*
g1877 not 1319(894) ; 1319(894)*
g1878 not 1320(904) ; 1320(904)*
g1879 not 1321(802) ; 1321(802)*
g1880 not 1322(809) ; 1322(809)*
g1881 not 1323(815) ; 1323(815)*
g1882 not 1299(825) ; 1299(825)*
g1883 not 1300(883) ; 1300(883)*
g1884 not 1301(893) ; 1301(893)*
g1885 not 1302(903) ; 1302(903)*
g1886 not 1303(803) ; 1303(803)*
g1887 not 1304(810) ; 1304(810)*
g1888 not 1305(816) ; 1305(816)*
g1889 not 1306(821) ; 1306(821)*
g1890 not 1282(829) ; 1282(829)*
g1891 not 1283(892) ; 1283(892)*
g1892 not 1284(902) ; 1284(902)*
g1893 not 1285(804) ; 1285(804)*
g1894 not 1286(811) ; 1286(811)*
g1895 not 1287(817) ; 1287(817)*
g1896 not 1288(822) ; 1288(822)*
g1897 not 1289(826) ; 1289(826)*
g1898 not 1265(832) ; 1265(832)*
g1899 not 1266(901) ; 1266(901)*
g1900 not 1267(805) ; 1267(805)*
g1901 not 1268(812) ; 1268(812)*
g1902 not 1269(818) ; 1269(818)*
g1903 not 1270(823) ; 1270(823)*
g1904 not 1271(827) ; 1271(827)*
g1905 not 1272(830) ; 1272(830)*
g1906 not 1248(834) ; 1248(834)*
g1907 not 1249(806) ; 1249(806)*
g1908 not 1250(813) ; 1250(813)*
g1909 not 1251(819) ; 1251(819)*
g1910 not 1252(824) ; 1252(824)*
g1911 not 1253(828) ; 1253(828)*
g1912 not 1254(831) ; 1254(831)*
g1913 not 1255(833) ; 1255(833)*
g1914 not 983(908) ; 983(908)*
g1915 not 984(408) ; 984(408)*
g1916 not 985(378) ; 985(378)*
g1917 not 1011(909) ; 1011(909)*
g1918 not 1012(386) ; 1012(386)*
g1919 not 1013(403) ; 1013(403)*
g1920 not 614(968) ; 614(968)*
g1921 not 616(424) ; 616(424)*
g1922 not 617(536) ; 617(536)*
g1923 not 2482(949) ; 2482(949)*
g1924 not 2483(999) ; 2483(999)*
g1925 not 2248(1006) ; 2248(1006)*
g1926 not 2251(1000) ; 2251(1000)*
g1927 not 2196(1007) ; 2196(1007)*
g1928 not 2199(1001) ; 2199(1001)*
g1929 not 2091(1008) ; 2091(1008)*
g1930 not 2094(1002) ; 2094(1002)*
g1931 not 2034(1009) ; 2034(1009)*
g1932 not 2037(1003) ; 2037(1003)*
g1933 not 1984(1010) ; 1984(1010)*
g1934 not 1987(1004) ; 1987(1004)*
g1935 not 1883(1011) ; 1883(1011)*
g1936 not 1886(1005) ; 1886(1005)*
g1937 not 2254(993) ; 2254(993)*
g1938 not 2255(987) ; 2255(987)*
g1939 not 2256(959) ; 2256(959)*
g1940 not 2202(994) ; 2202(994)*
g1941 not 2203(988) ; 2203(988)*
g1942 not 2204(961) ; 2204(961)*
g1943 not 2111(1035) ; 2111(1035)*
g1944 not 2114(388) ; 2114(388)*
g1945 not 2117(531) ; 2117(531)*
g1946 not 2097(995) ; 2097(995)*
g1947 not 2098(989) ; 2098(989)*
g1948 not 2099(963) ; 2099(963)*
g1949 not 2040(996) ; 2040(996)*
g1950 not 2041(990) ; 2041(990)*
g1951 not 2042(964) ; 2042(964)*
g1952 not 1990(997) ; 1990(997)*
g1953 not 1991(991) ; 1991(991)*
g1954 not 1992(966) ; 1992(966)*
g1955 not 1903(1034) ; 1903(1034)*
g1956 not 1906(411) ; 1906(411)*
g1957 not 1909(545) ; 1909(545)*
g1958 not 1889(998) ; 1889(998)*
g1959 not 1890(992) ; 1890(992)*
g1960 not 1891(967) ; 1891(967)*
g1961 not 1536(1016) ; 1536(1016)*
g1962 not 1537(1018) ; 1537(1018)*
g1963 not 1538(548) ; 1538(548)*
g1964 not 679(1015) ; 679(1015)*
g1965 not 680(420) ; 680(420)*
g1966 not 669(1019) ; 669(1019)*
g1967 not 671(426) ; 671(426)*
g1968 not 672(533) ; 672(533)*
g1969 not 1582(1020) ; 1582(1020)*
g1970 not 1583(1021) ; 1583(1021)*
g1971 not 1586(1022) ; 1586(1022)*
g1972 not 1587(1023) ; 1587(1023)*
g1973 not 1590(1024) ; 1590(1024)*
g1974 not 1591(1025) ; 1591(1025)*
g1975 not 1594(1026) ; 1594(1026)*
g1976 not 1595(1027) ; 1595(1027)*
g1977 not 1598(1028) ; 1598(1028)*
g1978 not 1599(1029) ; 1599(1029)*
g1979 not 1602(1030) ; 1602(1030)*
g1980 not 1603(1031) ; 1603(1031)*
g1981 not 1606(1032) ; 1606(1032)*
g1982 not 1607(1033) ; 1607(1033)*
g1983 not 661(1080) ; 661(1080)*
g1984 not 662(550) ; 662(550)*
g1985 not 2149(1104) ; 2149(1104)*
g1986 not 2150(1102) ; 2150(1102)*
g1987 not 2151(1122) ; 2151(1122)*
g1988 not 1939(1105) ; 1939(1105)*
g1989 not 1940(1103) ; 1940(1103)*
g1990 not 1941(1123) ; 1941(1123)*
g1991 not 2143(1116) ; 2143(1116)*
g1992 not 2146(1108) ; 2146(1108)*
g1993 not 1933(1117) ; 1933(1117)*
g1994 not 1936(1113) ; 1936(1113)*
g1995 not 689(1125) ; 689(1125)*
g1996 not 690(535) ; 690(535)*
g1997 not 691(524) ; 691(524)*
g1998 not 700(1160) ; 700(1160)*
g1999 not 701(523) ; 701(523)*
g2000 not 702(530) ; 702(530)*
g2001 not 2489(1100) ; 2489(1100)*
g2002 not 2490(1230) ; 2490(1230)*
g2003 not 2455(1095) ; 2455(1095)*
g2004 not 2518(1274) ; 2518(1274)*
g2005 not 2448(1099) ; 2448(1099)*
g2006 not 2517(1302) ; 2517(1302)*
g2007 not 2275(1246) ; 2275(1246)*
g2008 not 2500(1319) ; 2500(1319)*
g2009 not 1639(1130) ; 1639(1130)*
g2010 not 1641(1327) ; 1641(1327)*
g2011 not 1643(727) ; 1643(727)*
g2012 not 1630(1129) ; 1630(1129)*
g2013 not 1632(1326) ; 1632(1326)*
g2014 not 1634(730) ; 1634(730)*
g2015 not 1612(1127) ; 1612(1127)*
g2016 not 1614(1325) ; 1614(1325)*
g2017 not 1616(733) ; 1616(733)*
g2018 not 1648(1131) ; 1648(1131)*
g2019 not 1650(1322) ; 1650(1322)*
g2020 not 1652(1090) ; 1652(1090)*
g2021 not 1666(1133) ; 1666(1133)*
g2022 not 1668(1323) ; 1668(1323)*
g2023 not 1670(1225) ; 1670(1225)*
g2024 not 1675(1134) ; 1675(1134)*
g2025 not 1677(1324) ; 1677(1324)*
g2026 not 1679(1188) ; 1679(1188)*
g2027 not 2643(1328) ; 2643(1328)*
g2028 not 2645(1305) ; 2645(1305)*
g2029 not 1621(1128) ; 1621(1128)*
g2030 not 1623(1387) ; 1623(1387)*
g2031 not 1625(732) ; 1625(732)*
g2032 not 1657(1132) ; 1657(1132)*
g2033 not 1659(1386) ; 1659(1386)*
g2034 not 1661(1126) ; 1661(1126)*
g2035 not 397(1394) ; 397(1394)*
g2036 not 398(1366) ; 398(1366)*
g2037 not 929(734) ; 929(734)*
g2038 not 933(1419) ; 933(1419)*
g2039 not 938(722) ; 938(722)*
g2040 not 2633(1420) ; 2633(1420)*
g2041 not 2634(1416) ; 2634(1416)*
g2042 not 2805(1446) ; 2805(1446)*
g2043 not 2808(1443) ; 2808(1443)*
g2044 not 2811(1393) ; 2811(1393)*
g2045 not 2736(1502) ; 2736(1502)*
g2046 not 2739(1501) ; 2739(1501)*
g2047 not 2742(1390) ; 2742(1390)*
g2048 not 2600(1542) ; 2600(1542)*
g2049 not 2650(1404) ; 2650(1404)*
g2050 not 2661(1561) ; 2661(1561)*
g2051 not 2662(1548) ; 2662(1548)*
g2052 not 944(969) ; 944(969)*
g2053 not 947(910) ; 947(910)*
g2054 not 951(1564) ; 951(1564)*
g2055 not 2555(1566) ; 2555(1566)*
g2056 not 2638(1483) ; 2638(1483)*
g2057 not 2771(1523) ; 2771(1523)*
g2058 not 2774(1572) ; 2774(1572)*
g2059 not 2777(1445) ; 2777(1445)*
g2060 not 2788(1503) ; 2788(1503)*
g2061 not 2791(1573) ; 2791(1573)*
g2062 not 2794(1392) ; 2794(1392)*
g2063 not 2658(1575) ; 2658(1575)*
g2064 not 2659(1568) ; 2659(1568)*
g2065 not 2700(1520) ; 2700(1520)*
g2066 not 2703(1578) ; 2703(1578)*
g2067 not 2706(1444) ; 2706(1444)*
g2068 not 2754(1556) ; 2754(1556)*
g2069 not 2757(1579) ; 2757(1579)*
g2070 not 2760(1391) ; 2760(1391)*
g2071 not 2719(1538) ; 2719(1538)*
g2072 not 2722(1586) ; 2722(1586)*
g2073 not 2725(1389) ; 2725(1389)*
g2074 not 2681(1574) ; 2681(1574)*
g2075 not 2684(1596) ; 2684(1596)*
g2076 not 2687(1388) ; 2687(1388)*
g2077 not 2928(1623) ; 2928(1623)*
g2078 not 2929(1644) ; 2929(1644)*
g2079 not 2906(1677) ; 2906(1677)*
g2080 not 2907(1683) ; 2907(1683)*
g2081 not 2908(1676) ; 2908(1676)*
g2082 not 2909(1684) ; 2909(1684)*
