name C6288.iscas
i 1GAT(0)
i 18GAT(1)
i 35GAT(2)
i 52GAT(3)
i 69GAT(4)
i 86GAT(5)
i 103GAT(6)
i 120GAT(7)
i 137GAT(8)
i 154GAT(9)
i 171GAT(10)
i 188GAT(11)
i 205GAT(12)
i 222GAT(13)
i 239GAT(14)
i 256GAT(15)
i 273GAT(16)
i 290GAT(17)
i 307GAT(18)
i 324GAT(19)
i 341GAT(20)
i 358GAT(21)
i 375GAT(22)
i 392GAT(23)
i 409GAT(24)
i 426GAT(25)
i 443GAT(26)
i 460GAT(27)
i 477GAT(28)
i 494GAT(29)
i 511GAT(30)
i 528GAT(31)

o 545GAT(287)
o 1581GAT(423)
o 1901GAT(561)
o 2223GAT(700)
o 2548GAT(840)
o 2877GAT(983)
o 3211GAT(1128)
o 3552GAT(1275)
o 3895GAT(1423)
o 4241GAT(1572)
o 4591GAT(1722)
o 4946GAT(1876)
o 5308GAT(2031)
o 5672GAT(2187)
o 5971GAT(2309)
o 6123GAT(2368)
o 6150GAT(2378)
o 6160GAT(2383)
o 6170GAT(2388)
o 6180GAT(2393)
o 6190GAT(2398)
o 6200GAT(2403)
o 6210GAT(2408)
o 6220GAT(2413)
o 6230GAT(2418)
o 6240GAT(2423)
o 6250GAT(2428)
o 6260GAT(2433)
o 6270GAT(2438)
o 6280GAT(2443)
o 6287GAT(2444)
o 6288GAT(2447)

g1 and 528GAT(31) 256GAT(15) ; 1308GAT(32)
g2 and 511GAT(30) 256GAT(15) ; 1305GAT(33)
g3 and 494GAT(29) 256GAT(15) ; 1302GAT(34)
g4 and 477GAT(28) 256GAT(15) ; 1299GAT(35)
g5 and 460GAT(27) 256GAT(15) ; 1296GAT(36)
g6 and 443GAT(26) 256GAT(15) ; 1293GAT(37)
g7 and 426GAT(25) 256GAT(15) ; 1290GAT(38)
g8 and 409GAT(24) 256GAT(15) ; 1287GAT(39)
g9 and 392GAT(23) 256GAT(15) ; 1284GAT(40)
g10 and 375GAT(22) 256GAT(15) ; 1281GAT(41)
g11 and 358GAT(21) 256GAT(15) ; 1278GAT(42)
g12 and 341GAT(20) 256GAT(15) ; 1275GAT(43)
g13 and 324GAT(19) 256GAT(15) ; 1272GAT(44)
g14 and 307GAT(18) 256GAT(15) ; 1269GAT(45)
g15 and 290GAT(17) 256GAT(15) ; 1266GAT(46)
g16 and 273GAT(16) 256GAT(15) ; 1263GAT(47)
g17 and 528GAT(31) 239GAT(14) ; 1260GAT(48)
g18 and 511GAT(30) 239GAT(14) ; 1257GAT(49)
g19 and 494GAT(29) 239GAT(14) ; 1254GAT(50)
g20 and 477GAT(28) 239GAT(14) ; 1251GAT(51)
g21 and 460GAT(27) 239GAT(14) ; 1248GAT(52)
g22 and 443GAT(26) 239GAT(14) ; 1245GAT(53)
g23 and 426GAT(25) 239GAT(14) ; 1242GAT(54)
g24 and 409GAT(24) 239GAT(14) ; 1239GAT(55)
g25 and 392GAT(23) 239GAT(14) ; 1236GAT(56)
g26 and 375GAT(22) 239GAT(14) ; 1233GAT(57)
g27 and 358GAT(21) 239GAT(14) ; 1230GAT(58)
g28 and 341GAT(20) 239GAT(14) ; 1227GAT(59)
g29 and 324GAT(19) 239GAT(14) ; 1224GAT(60)
g30 and 307GAT(18) 239GAT(14) ; 1221GAT(61)
g31 and 290GAT(17) 239GAT(14) ; 1218GAT(62)
g32 and 273GAT(16) 239GAT(14) ; 1215GAT(63)
g33 and 528GAT(31) 222GAT(13) ; 1212GAT(64)
g34 and 511GAT(30) 222GAT(13) ; 1209GAT(65)
g35 and 494GAT(29) 222GAT(13) ; 1206GAT(66)
g36 and 477GAT(28) 222GAT(13) ; 1203GAT(67)
g37 and 460GAT(27) 222GAT(13) ; 1200GAT(68)
g38 and 443GAT(26) 222GAT(13) ; 1197GAT(69)
g39 and 426GAT(25) 222GAT(13) ; 1194GAT(70)
g40 and 409GAT(24) 222GAT(13) ; 1191GAT(71)
g41 and 392GAT(23) 222GAT(13) ; 1188GAT(72)
g42 and 375GAT(22) 222GAT(13) ; 1185GAT(73)
g43 and 358GAT(21) 222GAT(13) ; 1182GAT(74)
g44 and 341GAT(20) 222GAT(13) ; 1179GAT(75)
g45 and 324GAT(19) 222GAT(13) ; 1176GAT(76)
g46 and 307GAT(18) 222GAT(13) ; 1173GAT(77)
g47 and 290GAT(17) 222GAT(13) ; 1170GAT(78)
g48 and 273GAT(16) 222GAT(13) ; 1167GAT(79)
g49 and 528GAT(31) 205GAT(12) ; 1164GAT(80)
g50 and 511GAT(30) 205GAT(12) ; 1161GAT(81)
g51 and 494GAT(29) 205GAT(12) ; 1158GAT(82)
g52 and 477GAT(28) 205GAT(12) ; 1155GAT(83)
g53 and 460GAT(27) 205GAT(12) ; 1152GAT(84)
g54 and 443GAT(26) 205GAT(12) ; 1149GAT(85)
g55 and 426GAT(25) 205GAT(12) ; 1146GAT(86)
g56 and 409GAT(24) 205GAT(12) ; 1143GAT(87)
g57 and 392GAT(23) 205GAT(12) ; 1140GAT(88)
g58 and 375GAT(22) 205GAT(12) ; 1137GAT(89)
g59 and 358GAT(21) 205GAT(12) ; 1134GAT(90)
g60 and 341GAT(20) 205GAT(12) ; 1131GAT(91)
g61 and 324GAT(19) 205GAT(12) ; 1128GAT(92)
g62 and 307GAT(18) 205GAT(12) ; 1125GAT(93)
g63 and 290GAT(17) 205GAT(12) ; 1122GAT(94)
g64 and 273GAT(16) 205GAT(12) ; 1119GAT(95)
g65 and 528GAT(31) 188GAT(11) ; 1116GAT(96)
g66 and 511GAT(30) 188GAT(11) ; 1113GAT(97)
g67 and 494GAT(29) 188GAT(11) ; 1110GAT(98)
g68 and 477GAT(28) 188GAT(11) ; 1107GAT(99)
g69 and 460GAT(27) 188GAT(11) ; 1104GAT(100)
g70 and 443GAT(26) 188GAT(11) ; 1101GAT(101)
g71 and 426GAT(25) 188GAT(11) ; 1098GAT(102)
g72 and 409GAT(24) 188GAT(11) ; 1095GAT(103)
g73 and 392GAT(23) 188GAT(11) ; 1092GAT(104)
g74 and 375GAT(22) 188GAT(11) ; 1089GAT(105)
g75 and 358GAT(21) 188GAT(11) ; 1086GAT(106)
g76 and 341GAT(20) 188GAT(11) ; 1083GAT(107)
g77 and 324GAT(19) 188GAT(11) ; 1080GAT(108)
g78 and 307GAT(18) 188GAT(11) ; 1077GAT(109)
g79 and 290GAT(17) 188GAT(11) ; 1074GAT(110)
g80 and 273GAT(16) 188GAT(11) ; 1071GAT(111)
g81 and 528GAT(31) 171GAT(10) ; 1068GAT(112)
g82 and 511GAT(30) 171GAT(10) ; 1065GAT(113)
g83 and 494GAT(29) 171GAT(10) ; 1062GAT(114)
g84 and 477GAT(28) 171GAT(10) ; 1059GAT(115)
g85 and 460GAT(27) 171GAT(10) ; 1056GAT(116)
g86 and 443GAT(26) 171GAT(10) ; 1053GAT(117)
g87 and 426GAT(25) 171GAT(10) ; 1050GAT(118)
g88 and 409GAT(24) 171GAT(10) ; 1047GAT(119)
g89 and 392GAT(23) 171GAT(10) ; 1044GAT(120)
g90 and 375GAT(22) 171GAT(10) ; 1041GAT(121)
g91 and 358GAT(21) 171GAT(10) ; 1038GAT(122)
g92 and 341GAT(20) 171GAT(10) ; 1035GAT(123)
g93 and 324GAT(19) 171GAT(10) ; 1032GAT(124)
g94 and 307GAT(18) 171GAT(10) ; 1029GAT(125)
g95 and 290GAT(17) 171GAT(10) ; 1026GAT(126)
g96 and 273GAT(16) 171GAT(10) ; 1023GAT(127)
g97 and 528GAT(31) 154GAT(9) ; 1020GAT(128)
g98 and 511GAT(30) 154GAT(9) ; 1017GAT(129)
g99 and 494GAT(29) 154GAT(9) ; 1014GAT(130)
g100 and 477GAT(28) 154GAT(9) ; 1011GAT(131)
g101 and 460GAT(27) 154GAT(9) ; 1008GAT(132)
g102 and 443GAT(26) 154GAT(9) ; 1005GAT(133)
g103 and 426GAT(25) 154GAT(9) ; 1002GAT(134)
g104 and 409GAT(24) 154GAT(9) ; 999GAT(135)
g105 and 392GAT(23) 154GAT(9) ; 996GAT(136)
g106 and 375GAT(22) 154GAT(9) ; 993GAT(137)
g107 and 358GAT(21) 154GAT(9) ; 990GAT(138)
g108 and 341GAT(20) 154GAT(9) ; 987GAT(139)
g109 and 324GAT(19) 154GAT(9) ; 984GAT(140)
g110 and 307GAT(18) 154GAT(9) ; 981GAT(141)
g111 and 290GAT(17) 154GAT(9) ; 978GAT(142)
g112 and 273GAT(16) 154GAT(9) ; 975GAT(143)
g113 and 528GAT(31) 137GAT(8) ; 972GAT(144)
g114 and 511GAT(30) 137GAT(8) ; 969GAT(145)
g115 and 494GAT(29) 137GAT(8) ; 966GAT(146)
g116 and 477GAT(28) 137GAT(8) ; 963GAT(147)
g117 and 460GAT(27) 137GAT(8) ; 960GAT(148)
g118 and 443GAT(26) 137GAT(8) ; 957GAT(149)
g119 and 426GAT(25) 137GAT(8) ; 954GAT(150)
g120 and 409GAT(24) 137GAT(8) ; 951GAT(151)
g121 and 392GAT(23) 137GAT(8) ; 948GAT(152)
g122 and 375GAT(22) 137GAT(8) ; 945GAT(153)
g123 and 358GAT(21) 137GAT(8) ; 942GAT(154)
g124 and 341GAT(20) 137GAT(8) ; 939GAT(155)
g125 and 324GAT(19) 137GAT(8) ; 936GAT(156)
g126 and 307GAT(18) 137GAT(8) ; 933GAT(157)
g127 and 290GAT(17) 137GAT(8) ; 930GAT(158)
g128 and 273GAT(16) 137GAT(8) ; 927GAT(159)
g129 and 528GAT(31) 120GAT(7) ; 924GAT(160)
g130 and 511GAT(30) 120GAT(7) ; 921GAT(161)
g131 and 494GAT(29) 120GAT(7) ; 918GAT(162)
g132 and 477GAT(28) 120GAT(7) ; 915GAT(163)
g133 and 460GAT(27) 120GAT(7) ; 912GAT(164)
g134 and 443GAT(26) 120GAT(7) ; 909GAT(165)
g135 and 426GAT(25) 120GAT(7) ; 906GAT(166)
g136 and 409GAT(24) 120GAT(7) ; 903GAT(167)
g137 and 392GAT(23) 120GAT(7) ; 900GAT(168)
g138 and 375GAT(22) 120GAT(7) ; 897GAT(169)
g139 and 358GAT(21) 120GAT(7) ; 894GAT(170)
g140 and 341GAT(20) 120GAT(7) ; 891GAT(171)
g141 and 324GAT(19) 120GAT(7) ; 888GAT(172)
g142 and 307GAT(18) 120GAT(7) ; 885GAT(173)
g143 and 290GAT(17) 120GAT(7) ; 882GAT(174)
g144 and 273GAT(16) 120GAT(7) ; 879GAT(175)
g145 and 528GAT(31) 103GAT(6) ; 876GAT(176)
g146 and 511GAT(30) 103GAT(6) ; 873GAT(177)
g147 and 494GAT(29) 103GAT(6) ; 870GAT(178)
g148 and 477GAT(28) 103GAT(6) ; 867GAT(179)
g149 and 460GAT(27) 103GAT(6) ; 864GAT(180)
g150 and 443GAT(26) 103GAT(6) ; 861GAT(181)
g151 and 426GAT(25) 103GAT(6) ; 858GAT(182)
g152 and 409GAT(24) 103GAT(6) ; 855GAT(183)
g153 and 392GAT(23) 103GAT(6) ; 852GAT(184)
g154 and 375GAT(22) 103GAT(6) ; 849GAT(185)
g155 and 358GAT(21) 103GAT(6) ; 846GAT(186)
g156 and 341GAT(20) 103GAT(6) ; 843GAT(187)
g157 and 324GAT(19) 103GAT(6) ; 840GAT(188)
g158 and 307GAT(18) 103GAT(6) ; 837GAT(189)
g159 and 290GAT(17) 103GAT(6) ; 834GAT(190)
g160 and 273GAT(16) 103GAT(6) ; 831GAT(191)
g161 and 528GAT(31) 86GAT(5) ; 828GAT(192)
g162 and 511GAT(30) 86GAT(5) ; 825GAT(193)
g163 and 494GAT(29) 86GAT(5) ; 822GAT(194)
g164 and 477GAT(28) 86GAT(5) ; 819GAT(195)
g165 and 460GAT(27) 86GAT(5) ; 816GAT(196)
g166 and 443GAT(26) 86GAT(5) ; 813GAT(197)
g167 and 426GAT(25) 86GAT(5) ; 810GAT(198)
g168 and 409GAT(24) 86GAT(5) ; 807GAT(199)
g169 and 392GAT(23) 86GAT(5) ; 804GAT(200)
g170 and 375GAT(22) 86GAT(5) ; 801GAT(201)
g171 and 358GAT(21) 86GAT(5) ; 798GAT(202)
g172 and 341GAT(20) 86GAT(5) ; 795GAT(203)
g173 and 324GAT(19) 86GAT(5) ; 792GAT(204)
g174 and 307GAT(18) 86GAT(5) ; 789GAT(205)
g175 and 290GAT(17) 86GAT(5) ; 786GAT(206)
g176 and 273GAT(16) 86GAT(5) ; 783GAT(207)
g177 and 528GAT(31) 69GAT(4) ; 780GAT(208)
g178 and 511GAT(30) 69GAT(4) ; 777GAT(209)
g179 and 494GAT(29) 69GAT(4) ; 774GAT(210)
g180 and 477GAT(28) 69GAT(4) ; 771GAT(211)
g181 and 460GAT(27) 69GAT(4) ; 768GAT(212)
g182 and 443GAT(26) 69GAT(4) ; 765GAT(213)
g183 and 426GAT(25) 69GAT(4) ; 762GAT(214)
g184 and 409GAT(24) 69GAT(4) ; 759GAT(215)
g185 and 392GAT(23) 69GAT(4) ; 756GAT(216)
g186 and 375GAT(22) 69GAT(4) ; 753GAT(217)
g187 and 358GAT(21) 69GAT(4) ; 750GAT(218)
g188 and 341GAT(20) 69GAT(4) ; 747GAT(219)
g189 and 324GAT(19) 69GAT(4) ; 744GAT(220)
g190 and 307GAT(18) 69GAT(4) ; 741GAT(221)
g191 and 290GAT(17) 69GAT(4) ; 738GAT(222)
g192 and 273GAT(16) 69GAT(4) ; 735GAT(223)
g193 and 528GAT(31) 52GAT(3) ; 732GAT(224)
g194 and 511GAT(30) 52GAT(3) ; 729GAT(225)
g195 and 494GAT(29) 52GAT(3) ; 726GAT(226)
g196 and 477GAT(28) 52GAT(3) ; 723GAT(227)
g197 and 460GAT(27) 52GAT(3) ; 720GAT(228)
g198 and 443GAT(26) 52GAT(3) ; 717GAT(229)
g199 and 426GAT(25) 52GAT(3) ; 714GAT(230)
g200 and 409GAT(24) 52GAT(3) ; 711GAT(231)
g201 and 392GAT(23) 52GAT(3) ; 708GAT(232)
g202 and 375GAT(22) 52GAT(3) ; 705GAT(233)
g203 and 358GAT(21) 52GAT(3) ; 702GAT(234)
g204 and 341GAT(20) 52GAT(3) ; 699GAT(235)
g205 and 324GAT(19) 52GAT(3) ; 696GAT(236)
g206 and 307GAT(18) 52GAT(3) ; 693GAT(237)
g207 and 290GAT(17) 52GAT(3) ; 690GAT(238)
g208 and 273GAT(16) 52GAT(3) ; 687GAT(239)
g209 and 528GAT(31) 35GAT(2) ; 684GAT(240)
g210 and 511GAT(30) 35GAT(2) ; 681GAT(241)
g211 and 494GAT(29) 35GAT(2) ; 678GAT(242)
g212 and 477GAT(28) 35GAT(2) ; 675GAT(243)
g213 and 460GAT(27) 35GAT(2) ; 672GAT(244)
g214 and 443GAT(26) 35GAT(2) ; 669GAT(245)
g215 and 426GAT(25) 35GAT(2) ; 666GAT(246)
g216 and 409GAT(24) 35GAT(2) ; 663GAT(247)
g217 and 392GAT(23) 35GAT(2) ; 660GAT(248)
g218 and 375GAT(22) 35GAT(2) ; 657GAT(249)
g219 and 358GAT(21) 35GAT(2) ; 654GAT(250)
g220 and 341GAT(20) 35GAT(2) ; 651GAT(251)
g221 and 324GAT(19) 35GAT(2) ; 648GAT(252)
g222 and 307GAT(18) 35GAT(2) ; 645GAT(253)
g223 and 290GAT(17) 35GAT(2) ; 642GAT(254)
g224 and 273GAT(16) 35GAT(2) ; 639GAT(255)
g225 and 528GAT(31) 18GAT(1) ; 636GAT(256)
g226 and 511GAT(30) 18GAT(1) ; 633GAT(257)
g227 and 494GAT(29) 18GAT(1) ; 630GAT(258)
g228 and 477GAT(28) 18GAT(1) ; 627GAT(259)
g229 and 460GAT(27) 18GAT(1) ; 624GAT(260)
g230 and 443GAT(26) 18GAT(1) ; 621GAT(261)
g231 and 426GAT(25) 18GAT(1) ; 618GAT(262)
g232 and 409GAT(24) 18GAT(1) ; 615GAT(263)
g233 and 392GAT(23) 18GAT(1) ; 612GAT(264)
g234 and 375GAT(22) 18GAT(1) ; 609GAT(265)
g235 and 358GAT(21) 18GAT(1) ; 606GAT(266)
g236 and 341GAT(20) 18GAT(1) ; 603GAT(267)
g237 and 324GAT(19) 18GAT(1) ; 600GAT(268)
g238 and 307GAT(18) 18GAT(1) ; 597GAT(269)
g239 and 290GAT(17) 18GAT(1) ; 594GAT(270)
g240 and 273GAT(16) 18GAT(1) ; 591GAT(271)
g241 and 528GAT(31) 1GAT(0) ; 588GAT(272)
g242 and 511GAT(30) 1GAT(0) ; 585GAT(273)
g243 and 494GAT(29) 1GAT(0) ; 582GAT(274)
g244 and 477GAT(28) 1GAT(0) ; 579GAT(275)
g245 and 460GAT(27) 1GAT(0) ; 576GAT(276)
g246 and 443GAT(26) 1GAT(0) ; 573GAT(277)
g247 and 426GAT(25) 1GAT(0) ; 570GAT(278)
g248 and 409GAT(24) 1GAT(0) ; 567GAT(279)
g249 and 392GAT(23) 1GAT(0) ; 564GAT(280)
g250 and 375GAT(22) 1GAT(0) ; 561GAT(281)
g251 and 358GAT(21) 1GAT(0) ; 558GAT(282)
g252 and 341GAT(20) 1GAT(0) ; 555GAT(283)
g253 and 324GAT(19) 1GAT(0) ; 552GAT(284)
g254 and 307GAT(18) 1GAT(0) ; 549GAT(285)
g255 and 290GAT(17) 1GAT(0) ; 546GAT(286)
g256 and 273GAT(16) 1GAT(0) ; 545GAT(287)
g257 and 1263GAT(47) ; 1367GAT(288)
g258 and 1215GAT(63) ; 1363GAT(289)
g259 and 1167GAT(79) ; 1359GAT(290)
g260 and 1119GAT(95) ; 1355GAT(291)
g261 and 1071GAT(111) ; 1351GAT(292)
g262 and 1023GAT(127) ; 1347GAT(293)
g263 and 975GAT(143) ; 1343GAT(294)
g264 and 927GAT(159) ; 1339GAT(295)
g265 and 879GAT(175) ; 1335GAT(296)
g266 and 831GAT(191) ; 1331GAT(297)
g267 and 783GAT(207) ; 1327GAT(298)
g268 and 735GAT(223) ; 1323GAT(299)
g269 and 687GAT(239) ; 1319GAT(300)
g270 and 639GAT(255) ; 1315GAT(301)
g271 and 591GAT(271) ; 1311GAT(302)
g272 and 1367GAT(288) ; 1400GAT(303)
g273 and 1367GAT(288)* 1263GAT(47)* ; 1399GAT(304)
g274 and 1363GAT(289) ; 1398GAT(305)
g275 and 1363GAT(289)* 1215GAT(63)* ; 1397GAT(306)
g276 and 1359GAT(290) ; 1396GAT(307)
g277 and 1359GAT(290)* 1167GAT(79)* ; 1395GAT(308)
g278 and 1355GAT(291) ; 1394GAT(309)
g279 and 1355GAT(291)* 1119GAT(95)* ; 1393GAT(310)
g280 and 1351GAT(292) ; 1392GAT(311)
g281 and 1351GAT(292)* 1071GAT(111)* ; 1391GAT(312)
g282 and 1347GAT(293) ; 1390GAT(313)
g283 and 1347GAT(293)* 1023GAT(127)* ; 1389GAT(314)
g284 and 1343GAT(294) ; 1388GAT(315)
g285 and 1343GAT(294)* 975GAT(143)* ; 1387GAT(316)
g286 and 1339GAT(295) ; 1386GAT(317)
g287 and 1339GAT(295)* 927GAT(159)* ; 1385GAT(318)
g288 and 1335GAT(296) ; 1384GAT(319)
g289 and 1335GAT(296)* 879GAT(175)* ; 1383GAT(320)
g290 and 1331GAT(297) ; 1382GAT(321)
g291 and 1331GAT(297)* 831GAT(191)* ; 1381GAT(322)
g292 and 1327GAT(298) ; 1380GAT(323)
g293 and 1327GAT(298)* 783GAT(207)* ; 1379GAT(324)
g294 and 1323GAT(299) ; 1378GAT(325)
g295 and 1323GAT(299)* 735GAT(223)* ; 1377GAT(326)
g296 and 1319GAT(300) ; 1376GAT(327)
g297 and 1319GAT(300)* 687GAT(239)* ; 1375GAT(328)
g298 and 1315GAT(301) ; 1374GAT(329)
g299 and 1315GAT(301)* 639GAT(255)* ; 1373GAT(330)
g300 and 1311GAT(302) ; 1372GAT(331)
g301 and 1311GAT(302)* 591GAT(271)* ; 1371GAT(332)
g302 and 1400GAT(303)* 1399GAT(304)* ; 1443GAT(333)
g303 and 1398GAT(305)* 1397GAT(306)* ; 1440GAT(334)
g304 and 1396GAT(307)* 1395GAT(308)* ; 1437GAT(335)
g305 and 1394GAT(309)* 1393GAT(310)* ; 1434GAT(336)
g306 and 1392GAT(311)* 1391GAT(312)* ; 1431GAT(337)
g307 and 1390GAT(313)* 1389GAT(314)* ; 1428GAT(338)
g308 and 1388GAT(315)* 1387GAT(316)* ; 1425GAT(339)
g309 and 1386GAT(317)* 1385GAT(318)* ; 1422GAT(340)
g310 and 1384GAT(319)* 1383GAT(320)* ; 1419GAT(341)
g311 and 1382GAT(321)* 1381GAT(322)* ; 1416GAT(342)
g312 and 1380GAT(323)* 1379GAT(324)* ; 1413GAT(343)
g313 and 1378GAT(325)* 1377GAT(326)* ; 1410GAT(344)
g314 and 1376GAT(327)* 1375GAT(328)* ; 1407GAT(345)
g315 and 1374GAT(329)* 1373GAT(330)* ; 1404GAT(346)
g316 and 1372GAT(331)* 1371GAT(332)* ; 1401GAT(347)
g317 and 1218GAT(62)* 1443GAT(333)* ; 1502GAT(348)
g318 and 1170GAT(78)* 1440GAT(334)* ; 1498GAT(349)
g319 and 1122GAT(94)* 1437GAT(335)* ; 1494GAT(350)
g320 and 1074GAT(110)* 1434GAT(336)* ; 1490GAT(351)
g321 and 1026GAT(126)* 1431GAT(337)* ; 1486GAT(352)
g322 and 978GAT(142)* 1428GAT(338)* ; 1482GAT(353)
g323 and 930GAT(158)* 1425GAT(339)* ; 1478GAT(354)
g324 and 882GAT(174)* 1422GAT(340)* ; 1474GAT(355)
g325 and 834GAT(190)* 1419GAT(341)* ; 1470GAT(356)
g326 and 786GAT(206)* 1416GAT(342)* ; 1466GAT(357)
g327 and 738GAT(222)* 1413GAT(343)* ; 1462GAT(358)
g328 and 690GAT(238)* 1410GAT(344)* ; 1458GAT(359)
g329 and 642GAT(254)* 1407GAT(345)* ; 1454GAT(360)
g330 and 594GAT(270)* 1404GAT(346)* ; 1450GAT(361)
g331 and 546GAT(286)* 1401GAT(347)* ; 1446GAT(362)
g332 and 1502GAT(348)* 1367GAT(288)* ; 1578GAT(363)
g333 and 1502GAT(348)* 1443GAT(333)* ; 1576GAT(364)
g334 and 1218GAT(62)* 1502GAT(348)* ; 1577GAT(365)
g335 and 1498GAT(349)* 1363GAT(289)* ; 1573GAT(366)
g336 and 1498GAT(349)* 1440GAT(334)* ; 1571GAT(367)
g337 and 1170GAT(78)* 1498GAT(349)* ; 1572GAT(368)
g338 and 1494GAT(350)* 1359GAT(290)* ; 1568GAT(369)
g339 and 1494GAT(350)* 1437GAT(335)* ; 1566GAT(370)
g340 and 1122GAT(94)* 1494GAT(350)* ; 1567GAT(371)
g341 and 1490GAT(351)* 1355GAT(291)* ; 1563GAT(372)
g342 and 1490GAT(351)* 1434GAT(336)* ; 1561GAT(373)
g343 and 1074GAT(110)* 1490GAT(351)* ; 1562GAT(374)
g344 and 1486GAT(352)* 1351GAT(292)* ; 1558GAT(375)
g345 and 1486GAT(352)* 1431GAT(337)* ; 1556GAT(376)
g346 and 1026GAT(126)* 1486GAT(352)* ; 1557GAT(377)
g347 and 1482GAT(353)* 1347GAT(293)* ; 1553GAT(378)
g348 and 1482GAT(353)* 1428GAT(338)* ; 1551GAT(379)
g349 and 978GAT(142)* 1482GAT(353)* ; 1552GAT(380)
g350 and 1478GAT(354)* 1343GAT(294)* ; 1548GAT(381)
g351 and 1478GAT(354)* 1425GAT(339)* ; 1546GAT(382)
g352 and 930GAT(158)* 1478GAT(354)* ; 1547GAT(383)
g353 and 1474GAT(355)* 1339GAT(295)* ; 1543GAT(384)
g354 and 1474GAT(355)* 1422GAT(340)* ; 1541GAT(385)
g355 and 882GAT(174)* 1474GAT(355)* ; 1542GAT(386)
g356 and 1470GAT(356)* 1335GAT(296)* ; 1538GAT(387)
g357 and 1470GAT(356)* 1419GAT(341)* ; 1536GAT(388)
g358 and 834GAT(190)* 1470GAT(356)* ; 1537GAT(389)
g359 and 1466GAT(357)* 1331GAT(297)* ; 1533GAT(390)
g360 and 1466GAT(357)* 1416GAT(342)* ; 1531GAT(391)
g361 and 786GAT(206)* 1466GAT(357)* ; 1532GAT(392)
g362 and 1462GAT(358)* 1327GAT(298)* ; 1528GAT(393)
g363 and 1462GAT(358)* 1413GAT(343)* ; 1526GAT(394)
g364 and 738GAT(222)* 1462GAT(358)* ; 1527GAT(395)
g365 and 1458GAT(359)* 1323GAT(299)* ; 1523GAT(396)
g366 and 1458GAT(359)* 1410GAT(344)* ; 1521GAT(397)
g367 and 690GAT(238)* 1458GAT(359)* ; 1522GAT(398)
g368 and 1454GAT(360)* 1319GAT(300)* ; 1518GAT(399)
g369 and 1454GAT(360)* 1407GAT(345)* ; 1516GAT(400)
g370 and 642GAT(254)* 1454GAT(360)* ; 1517GAT(401)
g371 and 1450GAT(361)* 1315GAT(301)* ; 1513GAT(402)
g372 and 1450GAT(361)* 1404GAT(346)* ; 1511GAT(403)
g373 and 594GAT(270)* 1450GAT(361)* ; 1512GAT(404)
g374 and 1446GAT(362)* 1311GAT(302)* ; 1508GAT(405)
g375 and 1446GAT(362)* 1401GAT(347)* ; 1506GAT(406)
g376 and 546GAT(286)* 1446GAT(362)* ; 1507GAT(407)
g377 and 1578GAT(363)* 1266GAT(46)* ; 1624GAT(408)
g378 and 1577GAT(365)* 1576GAT(364)* ; 1621GAT(409)
g379 and 1572GAT(368)* 1571GAT(367)* ; 1618GAT(410)
g380 and 1567GAT(371)* 1566GAT(370)* ; 1615GAT(411)
g381 and 1562GAT(374)* 1561GAT(373)* ; 1612GAT(412)
g382 and 1557GAT(377)* 1556GAT(376)* ; 1609GAT(413)
g383 and 1552GAT(380)* 1551GAT(379)* ; 1606GAT(414)
g384 and 1547GAT(383)* 1546GAT(382)* ; 1603GAT(415)
g385 and 1542GAT(386)* 1541GAT(385)* ; 1600GAT(416)
g386 and 1537GAT(389)* 1536GAT(388)* ; 1597GAT(417)
g387 and 1532GAT(392)* 1531GAT(391)* ; 1594GAT(418)
g388 and 1527GAT(395)* 1526GAT(394)* ; 1591GAT(419)
g389 and 1522GAT(398)* 1521GAT(397)* ; 1588GAT(420)
g390 and 1517GAT(401)* 1516GAT(400)* ; 1585GAT(421)
g391 and 1512GAT(404)* 1511GAT(403)* ; 1582GAT(422)
g392 and 1507GAT(407)* 1506GAT(406)* ; 1581GAT(423)
g393 and 1624GAT(408)* 1266GAT(46)* ; 1684GAT(424)
g394 and 1578GAT(363)* 1624GAT(408)* ; 1685GAT(425)
g395 and 1573GAT(366)* 1621GAT(409)* ; 1680GAT(426)
g396 and 1568GAT(369)* 1618GAT(410)* ; 1676GAT(427)
g397 and 1563GAT(372)* 1615GAT(411)* ; 1672GAT(428)
g398 and 1558GAT(375)* 1612GAT(412)* ; 1668GAT(429)
g399 and 1553GAT(378)* 1609GAT(413)* ; 1664GAT(430)
g400 and 1548GAT(381)* 1606GAT(414)* ; 1660GAT(431)
g401 and 1543GAT(384)* 1603GAT(415)* ; 1656GAT(432)
g402 and 1538GAT(387)* 1600GAT(416)* ; 1652GAT(433)
g403 and 1533GAT(390)* 1597GAT(417)* ; 1648GAT(434)
g404 and 1528GAT(393)* 1594GAT(418)* ; 1644GAT(435)
g405 and 1523GAT(396)* 1591GAT(419)* ; 1640GAT(436)
g406 and 1518GAT(399)* 1588GAT(420)* ; 1636GAT(437)
g407 and 1513GAT(402)* 1585GAT(421)* ; 1632GAT(438)
g408 and 1508GAT(405)* 1582GAT(422)* ; 1628GAT(439)
g409 and 1685GAT(425)* 1684GAT(424)* ; 1714GAT(440)
g410 and 1680GAT(426)* 1621GAT(409)* ; 1712GAT(441)
g411 and 1573GAT(366)* 1680GAT(426)* ; 1713GAT(442)
g412 and 1676GAT(427)* 1618GAT(410)* ; 1710GAT(443)
g413 and 1568GAT(369)* 1676GAT(427)* ; 1711GAT(444)
g414 and 1672GAT(428)* 1615GAT(411)* ; 1708GAT(445)
g415 and 1563GAT(372)* 1672GAT(428)* ; 1709GAT(446)
g416 and 1668GAT(429)* 1612GAT(412)* ; 1706GAT(447)
g417 and 1558GAT(375)* 1668GAT(429)* ; 1707GAT(448)
g418 and 1664GAT(430)* 1609GAT(413)* ; 1704GAT(449)
g419 and 1553GAT(378)* 1664GAT(430)* ; 1705GAT(450)
g420 and 1660GAT(431)* 1606GAT(414)* ; 1702GAT(451)
g421 and 1548GAT(381)* 1660GAT(431)* ; 1703GAT(452)
g422 and 1656GAT(432)* 1603GAT(415)* ; 1700GAT(453)
g423 and 1543GAT(384)* 1656GAT(432)* ; 1701GAT(454)
g424 and 1652GAT(433)* 1600GAT(416)* ; 1698GAT(455)
g425 and 1538GAT(387)* 1652GAT(433)* ; 1699GAT(456)
g426 and 1648GAT(434)* 1597GAT(417)* ; 1696GAT(457)
g427 and 1533GAT(390)* 1648GAT(434)* ; 1697GAT(458)
g428 and 1644GAT(435)* 1594GAT(418)* ; 1694GAT(459)
g429 and 1528GAT(393)* 1644GAT(435)* ; 1695GAT(460)
g430 and 1640GAT(436)* 1591GAT(419)* ; 1692GAT(461)
g431 and 1523GAT(396)* 1640GAT(436)* ; 1693GAT(462)
g432 and 1636GAT(437)* 1588GAT(420)* ; 1690GAT(463)
g433 and 1518GAT(399)* 1636GAT(437)* ; 1691GAT(464)
g434 and 1632GAT(438)* 1585GAT(421)* ; 1688GAT(465)
g435 and 1513GAT(402)* 1632GAT(438)* ; 1689GAT(466)
g436 and 1628GAT(439)* 1582GAT(422)* ; 1686GAT(467)
g437 and 1508GAT(405)* 1628GAT(439)* ; 1687GAT(468)
g438 and 1713GAT(442)* 1712GAT(441)* ; 1756GAT(469)
g439 and 1221GAT(61)* 1714GAT(440)* ; 1759GAT(470)
g440 and 1711GAT(444)* 1710GAT(443)* ; 1753GAT(471)
g441 and 1709GAT(446)* 1708GAT(445)* ; 1750GAT(472)
g442 and 1707GAT(448)* 1706GAT(447)* ; 1747GAT(473)
g443 and 1705GAT(450)* 1704GAT(449)* ; 1744GAT(474)
g444 and 1703GAT(452)* 1702GAT(451)* ; 1741GAT(475)
g445 and 1701GAT(454)* 1700GAT(453)* ; 1738GAT(476)
g446 and 1699GAT(456)* 1698GAT(455)* ; 1735GAT(477)
g447 and 1697GAT(458)* 1696GAT(457)* ; 1732GAT(478)
g448 and 1695GAT(460)* 1694GAT(459)* ; 1729GAT(479)
g449 and 1693GAT(462)* 1692GAT(461)* ; 1726GAT(480)
g450 and 1691GAT(464)* 1690GAT(463)* ; 1723GAT(481)
g451 and 1689GAT(466)* 1688GAT(465)* ; 1720GAT(482)
g452 and 1687GAT(468)* 1686GAT(467)* ; 1717GAT(483)
g453 and 1759GAT(470)* 1624GAT(408)* ; 1821GAT(484)
g454 and 1759GAT(470)* 1714GAT(440)* ; 1819GAT(485)
g455 and 1221GAT(61)* 1759GAT(470)* ; 1820GAT(486)
g456 and 1173GAT(77)* 1756GAT(469)* ; 1815GAT(487)
g457 and 1125GAT(93)* 1753GAT(471)* ; 1811GAT(488)
g458 and 1077GAT(109)* 1750GAT(472)* ; 1807GAT(489)
g459 and 1029GAT(125)* 1747GAT(473)* ; 1803GAT(490)
g460 and 981GAT(141)* 1744GAT(474)* ; 1799GAT(491)
g461 and 933GAT(157)* 1741GAT(475)* ; 1795GAT(492)
g462 and 885GAT(173)* 1738GAT(476)* ; 1791GAT(493)
g463 and 837GAT(189)* 1735GAT(477)* ; 1787GAT(494)
g464 and 789GAT(205)* 1732GAT(478)* ; 1783GAT(495)
g465 and 741GAT(221)* 1729GAT(479)* ; 1779GAT(496)
g466 and 693GAT(237)* 1726GAT(480)* ; 1775GAT(497)
g467 and 645GAT(253)* 1723GAT(481)* ; 1771GAT(498)
g468 and 597GAT(269)* 1720GAT(482)* ; 1767GAT(499)
g469 and 549GAT(285)* 1717GAT(483)* ; 1763GAT(500)
g470 and 1821GAT(484)* 1269GAT(45)* ; 1897GAT(501)
g471 and 1820GAT(486)* 1819GAT(485)* ; 1894GAT(502)
g472 and 1815GAT(487)* 1756GAT(469)* ; 1889GAT(503)
g473 and 1815GAT(487)* 1680GAT(426)* ; 1891GAT(504)
g474 and 1811GAT(488)* 1753GAT(471)* ; 1884GAT(505)
g475 and 1173GAT(77)* 1815GAT(487)* ; 1890GAT(506)
g476 and 1811GAT(488)* 1676GAT(427)* ; 1886GAT(507)
g477 and 1807GAT(489)* 1750GAT(472)* ; 1879GAT(508)
g478 and 1125GAT(93)* 1811GAT(488)* ; 1885GAT(509)
g479 and 1807GAT(489)* 1672GAT(428)* ; 1881GAT(510)
g480 and 1803GAT(490)* 1747GAT(473)* ; 1874GAT(511)
g481 and 1077GAT(109)* 1807GAT(489)* ; 1880GAT(512)
g482 and 1803GAT(490)* 1668GAT(429)* ; 1876GAT(513)
g483 and 1799GAT(491)* 1744GAT(474)* ; 1869GAT(514)
g484 and 1029GAT(125)* 1803GAT(490)* ; 1875GAT(515)
g485 and 1799GAT(491)* 1664GAT(430)* ; 1871GAT(516)
g486 and 1795GAT(492)* 1741GAT(475)* ; 1864GAT(517)
g487 and 981GAT(141)* 1799GAT(491)* ; 1870GAT(518)
g488 and 1795GAT(492)* 1660GAT(431)* ; 1866GAT(519)
g489 and 1791GAT(493)* 1738GAT(476)* ; 1859GAT(520)
g490 and 933GAT(157)* 1795GAT(492)* ; 1865GAT(521)
g491 and 1791GAT(493)* 1656GAT(432)* ; 1861GAT(522)
g492 and 1787GAT(494)* 1735GAT(477)* ; 1854GAT(523)
g493 and 885GAT(173)* 1791GAT(493)* ; 1860GAT(524)
g494 and 1787GAT(494)* 1652GAT(433)* ; 1856GAT(525)
g495 and 1783GAT(495)* 1732GAT(478)* ; 1849GAT(526)
g496 and 837GAT(189)* 1787GAT(494)* ; 1855GAT(527)
g497 and 1783GAT(495)* 1648GAT(434)* ; 1851GAT(528)
g498 and 1779GAT(496)* 1729GAT(479)* ; 1844GAT(529)
g499 and 789GAT(205)* 1783GAT(495)* ; 1850GAT(530)
g500 and 1779GAT(496)* 1644GAT(435)* ; 1846GAT(531)
g501 and 1775GAT(497)* 1726GAT(480)* ; 1839GAT(532)
g502 and 741GAT(221)* 1779GAT(496)* ; 1845GAT(533)
g503 and 1775GAT(497)* 1640GAT(436)* ; 1841GAT(534)
g504 and 1771GAT(498)* 1723GAT(481)* ; 1834GAT(535)
g505 and 693GAT(237)* 1775GAT(497)* ; 1840GAT(536)
g506 and 1771GAT(498)* 1636GAT(437)* ; 1836GAT(537)
g507 and 1767GAT(499)* 1720GAT(482)* ; 1829GAT(538)
g508 and 645GAT(253)* 1771GAT(498)* ; 1835GAT(539)
g509 and 1767GAT(499)* 1632GAT(438)* ; 1831GAT(540)
g510 and 1763GAT(500)* 1717GAT(483)* ; 1824GAT(541)
g511 and 597GAT(269)* 1767GAT(499)* ; 1830GAT(542)
g512 and 1763GAT(500)* 1628GAT(439)* ; 1826GAT(543)
g513 and 549GAT(285)* 1763GAT(500)* ; 1825GAT(544)
g514 and 1897GAT(501)* 1269GAT(45)* ; 1945GAT(545)
g515 and 1821GAT(484)* 1897GAT(501)* ; 1946GAT(546)
g516 and 1891GAT(504)* 1894GAT(502)* ; 1941GAT(547)
g517 and 1890GAT(506)* 1889GAT(503)* ; 1938GAT(548)
g518 and 1885GAT(509)* 1884GAT(505)* ; 1935GAT(549)
g519 and 1880GAT(512)* 1879GAT(508)* ; 1932GAT(550)
g520 and 1875GAT(515)* 1874GAT(511)* ; 1929GAT(551)
g521 and 1870GAT(518)* 1869GAT(514)* ; 1926GAT(552)
g522 and 1865GAT(521)* 1864GAT(517)* ; 1923GAT(553)
g523 and 1860GAT(524)* 1859GAT(520)* ; 1920GAT(554)
g524 and 1855GAT(527)* 1854GAT(523)* ; 1917GAT(555)
g525 and 1850GAT(530)* 1849GAT(526)* ; 1914GAT(556)
g526 and 1845GAT(533)* 1844GAT(529)* ; 1911GAT(557)
g527 and 1840GAT(536)* 1839GAT(532)* ; 1908GAT(558)
g528 and 1835GAT(539)* 1834GAT(535)* ; 1905GAT(559)
g529 and 1830GAT(542)* 1829GAT(538)* ; 1902GAT(560)
g530 and 1825GAT(544)* 1824GAT(541)* ; 1901GAT(561)
g531 and 1946GAT(546)* 1945GAT(545)* ; 2001GAT(562)
g532 and 1941GAT(547)* 1894GAT(502)* ; 1999GAT(563)
g533 and 1891GAT(504)* 1941GAT(547)* ; 2000GAT(564)
g534 and 1886GAT(507)* 1938GAT(548)* ; 1995GAT(565)
g535 and 1881GAT(510)* 1935GAT(549)* ; 1991GAT(566)
g536 and 1876GAT(513)* 1932GAT(550)* ; 1987GAT(567)
g537 and 1871GAT(516)* 1929GAT(551)* ; 1983GAT(568)
g538 and 1866GAT(519)* 1926GAT(552)* ; 1979GAT(569)
g539 and 1861GAT(522)* 1923GAT(553)* ; 1975GAT(570)
g540 and 1856GAT(525)* 1920GAT(554)* ; 1971GAT(571)
g541 and 1851GAT(528)* 1917GAT(555)* ; 1967GAT(572)
g542 and 1846GAT(531)* 1914GAT(556)* ; 1963GAT(573)
g543 and 1841GAT(534)* 1911GAT(557)* ; 1959GAT(574)
g544 and 1836GAT(537)* 1908GAT(558)* ; 1955GAT(575)
g545 and 1831GAT(540)* 1905GAT(559)* ; 1951GAT(576)
g546 and 1826GAT(543)* 1902GAT(560)* ; 1947GAT(577)
g547 and 2000GAT(564)* 1999GAT(563)* ; 2030GAT(578)
g548 and 1995GAT(565)* 1938GAT(548)* ; 2028GAT(579)
g549 and 1224GAT(60)* 2001GAT(562)* ; 2033GAT(580)
g550 and 1991GAT(566)* 1935GAT(549)* ; 2026GAT(581)
g551 and 1886GAT(507)* 1995GAT(565)* ; 2029GAT(582)
g552 and 1987GAT(567)* 1932GAT(550)* ; 2024GAT(583)
g553 and 1881GAT(510)* 1991GAT(566)* ; 2027GAT(584)
g554 and 1983GAT(568)* 1929GAT(551)* ; 2022GAT(585)
g555 and 1876GAT(513)* 1987GAT(567)* ; 2025GAT(586)
g556 and 1979GAT(569)* 1926GAT(552)* ; 2020GAT(587)
g557 and 1871GAT(516)* 1983GAT(568)* ; 2023GAT(588)
g558 and 1975GAT(570)* 1923GAT(553)* ; 2018GAT(589)
g559 and 1866GAT(519)* 1979GAT(569)* ; 2021GAT(590)
g560 and 1971GAT(571)* 1920GAT(554)* ; 2016GAT(591)
g561 and 1861GAT(522)* 1975GAT(570)* ; 2019GAT(592)
g562 and 1967GAT(572)* 1917GAT(555)* ; 2014GAT(593)
g563 and 1856GAT(525)* 1971GAT(571)* ; 2017GAT(594)
g564 and 1963GAT(573)* 1914GAT(556)* ; 2012GAT(595)
g565 and 1851GAT(528)* 1967GAT(572)* ; 2015GAT(596)
g566 and 1959GAT(574)* 1911GAT(557)* ; 2010GAT(597)
g567 and 1846GAT(531)* 1963GAT(573)* ; 2013GAT(598)
g568 and 1955GAT(575)* 1908GAT(558)* ; 2008GAT(599)
g569 and 1841GAT(534)* 1959GAT(574)* ; 2011GAT(600)
g570 and 1951GAT(576)* 1905GAT(559)* ; 2006GAT(601)
g571 and 1836GAT(537)* 1955GAT(575)* ; 2009GAT(602)
g572 and 1947GAT(577)* 1902GAT(560)* ; 2004GAT(603)
g573 and 1831GAT(540)* 1951GAT(576)* ; 2007GAT(604)
g574 and 1826GAT(543)* 1947GAT(577)* ; 2005GAT(605)
g575 and 2033GAT(580)* 1897GAT(501)* ; 2082GAT(606)
g576 and 2033GAT(580)* 2001GAT(562)* ; 2080GAT(607)
g577 and 2029GAT(582)* 2028GAT(579)* ; 2073GAT(608)
g578 and 1224GAT(60)* 2033GAT(580)* ; 2081GAT(609)
g579 and 2027GAT(584)* 2026GAT(581)* ; 2070GAT(610)
g580 and 1176GAT(76)* 2030GAT(578)* ; 2076GAT(611)
g581 and 2025GAT(586)* 2024GAT(583)* ; 2067GAT(612)
g582 and 2023GAT(588)* 2022GAT(585)* ; 2064GAT(613)
g583 and 2021GAT(590)* 2020GAT(587)* ; 2061GAT(614)
g584 and 2019GAT(592)* 2018GAT(589)* ; 2058GAT(615)
g585 and 2017GAT(594)* 2016GAT(591)* ; 2055GAT(616)
g586 and 2015GAT(596)* 2014GAT(593)* ; 2052GAT(617)
g587 and 2013GAT(598)* 2012GAT(595)* ; 2049GAT(618)
g588 and 2011GAT(600)* 2010GAT(597)* ; 2046GAT(619)
g589 and 2009GAT(602)* 2008GAT(599)* ; 2043GAT(620)
g590 and 2007GAT(604)* 2006GAT(601)* ; 2040GAT(621)
g591 and 2005GAT(605)* 2004GAT(603)* ; 2037GAT(622)
g592 and 2082GAT(606)* 1272GAT(44)* ; 2145GAT(623)
g593 and 2081GAT(609)* 2080GAT(607)* ; 2142GAT(624)
g594 and 2076GAT(611)* 1941GAT(547)* ; 2139GAT(625)
g595 and 2076GAT(611)* 2030GAT(578)* ; 2137GAT(626)
g596 and 1176GAT(76)* 2076GAT(611)* ; 2138GAT(627)
g597 and 1128GAT(92)* 2073GAT(608)* ; 2133GAT(628)
g598 and 1080GAT(108)* 2070GAT(610)* ; 2129GAT(629)
g599 and 1032GAT(124)* 2067GAT(612)* ; 2125GAT(630)
g600 and 984GAT(140)* 2064GAT(613)* ; 2121GAT(631)
g601 and 936GAT(156)* 2061GAT(614)* ; 2117GAT(632)
g602 and 888GAT(172)* 2058GAT(615)* ; 2113GAT(633)
g603 and 840GAT(188)* 2055GAT(616)* ; 2109GAT(634)
g604 and 792GAT(204)* 2052GAT(617)* ; 2105GAT(635)
g605 and 744GAT(220)* 2049GAT(618)* ; 2101GAT(636)
g606 and 696GAT(236)* 2046GAT(619)* ; 2097GAT(637)
g607 and 648GAT(252)* 2043GAT(620)* ; 2093GAT(638)
g608 and 600GAT(268)* 2040GAT(621)* ; 2089GAT(639)
g609 and 552GAT(284)* 2037GAT(622)* ; 2085GAT(640)
g610 and 2145GAT(623)* 1272GAT(44)* ; 2221GAT(641)
g611 and 2082GAT(606)* 2145GAT(623)* ; 2222GAT(642)
g612 and 2139GAT(625)* 2142GAT(624)* ; 2217GAT(643)
g613 and 2138GAT(627)* 2137GAT(626)* ; 2214GAT(644)
g614 and 2133GAT(628)* 2073GAT(608)* ; 2209GAT(645)
g615 and 2129GAT(629)* 2070GAT(610)* ; 2204GAT(646)
g616 and 2133GAT(628)* 1995GAT(565)* ; 2211GAT(647)
g617 and 2125GAT(630)* 2067GAT(612)* ; 2199GAT(648)
g618 and 1128GAT(92)* 2133GAT(628)* ; 2210GAT(649)
g619 and 2129GAT(629)* 1991GAT(566)* ; 2206GAT(650)
g620 and 2121GAT(631)* 2064GAT(613)* ; 2194GAT(651)
g621 and 1080GAT(108)* 2129GAT(629)* ; 2205GAT(652)
g622 and 2125GAT(630)* 1987GAT(567)* ; 2201GAT(653)
g623 and 2117GAT(632)* 2061GAT(614)* ; 2189GAT(654)
g624 and 1032GAT(124)* 2125GAT(630)* ; 2200GAT(655)
g625 and 2121GAT(631)* 1983GAT(568)* ; 2196GAT(656)
g626 and 2113GAT(633)* 2058GAT(615)* ; 2184GAT(657)
g627 and 984GAT(140)* 2121GAT(631)* ; 2195GAT(658)
g628 and 2117GAT(632)* 1979GAT(569)* ; 2191GAT(659)
g629 and 2109GAT(634)* 2055GAT(616)* ; 2179GAT(660)
g630 and 936GAT(156)* 2117GAT(632)* ; 2190GAT(661)
g631 and 2113GAT(633)* 1975GAT(570)* ; 2186GAT(662)
g632 and 2105GAT(635)* 2052GAT(617)* ; 2174GAT(663)
g633 and 888GAT(172)* 2113GAT(633)* ; 2185GAT(664)
g634 and 2109GAT(634)* 1971GAT(571)* ; 2181GAT(665)
g635 and 2101GAT(636)* 2049GAT(618)* ; 2169GAT(666)
g636 and 840GAT(188)* 2109GAT(634)* ; 2180GAT(667)
g637 and 2105GAT(635)* 1967GAT(572)* ; 2176GAT(668)
g638 and 2097GAT(637)* 2046GAT(619)* ; 2164GAT(669)
g639 and 792GAT(204)* 2105GAT(635)* ; 2175GAT(670)
g640 and 2101GAT(636)* 1963GAT(573)* ; 2171GAT(671)
g641 and 2093GAT(638)* 2043GAT(620)* ; 2159GAT(672)
g642 and 744GAT(220)* 2101GAT(636)* ; 2170GAT(673)
g643 and 2097GAT(637)* 1959GAT(574)* ; 2166GAT(674)
g644 and 2089GAT(639)* 2040GAT(621)* ; 2154GAT(675)
g645 and 696GAT(236)* 2097GAT(637)* ; 2165GAT(676)
g646 and 2093GAT(638)* 1955GAT(575)* ; 2161GAT(677)
g647 and 2085GAT(640)* 2037GAT(622)* ; 2149GAT(678)
g648 and 648GAT(252)* 2093GAT(638)* ; 2160GAT(679)
g649 and 2089GAT(639)* 1951GAT(576)* ; 2156GAT(680)
g650 and 600GAT(268)* 2089GAT(639)* ; 2155GAT(681)
g651 and 2085GAT(640)* 1947GAT(577)* ; 2151GAT(682)
g652 and 552GAT(284)* 2085GAT(640)* ; 2150GAT(683)
g653 and 2222GAT(642)* 2221GAT(641)* ; 2266GAT(684)
g654 and 2217GAT(643)* 2142GAT(624)* ; 2264GAT(685)
g655 and 2139GAT(625)* 2217GAT(643)* ; 2265GAT(686)
g656 and 2211GAT(647)* 2214GAT(644)* ; 2260GAT(687)
g657 and 2210GAT(649)* 2209GAT(645)* ; 2257GAT(688)
g658 and 2205GAT(652)* 2204GAT(646)* ; 2254GAT(689)
g659 and 2200GAT(655)* 2199GAT(648)* ; 2251GAT(690)
g660 and 2195GAT(658)* 2194GAT(651)* ; 2248GAT(691)
g661 and 2190GAT(661)* 2189GAT(654)* ; 2245GAT(692)
g662 and 2185GAT(664)* 2184GAT(657)* ; 2242GAT(693)
g663 and 2180GAT(667)* 2179GAT(660)* ; 2239GAT(694)
g664 and 2175GAT(670)* 2174GAT(663)* ; 2236GAT(695)
g665 and 2170GAT(673)* 2169GAT(666)* ; 2233GAT(696)
g666 and 2165GAT(676)* 2164GAT(669)* ; 2230GAT(697)
g667 and 2160GAT(679)* 2159GAT(672)* ; 2227GAT(698)
g668 and 2155GAT(681)* 2154GAT(675)* ; 2224GAT(699)
g669 and 2150GAT(683)* 2149GAT(678)* ; 2223GAT(700)
g670 and 2265GAT(686)* 2264GAT(685)* ; 2319GAT(701)
g671 and 2260GAT(687)* 2214GAT(644)* ; 2317GAT(702)
g672 and 1227GAT(59)* 2266GAT(684)* ; 2322GAT(703)
g673 and 2211GAT(647)* 2260GAT(687)* ; 2318GAT(704)
g674 and 2206GAT(650)* 2257GAT(688)* ; 2313GAT(705)
g675 and 2201GAT(653)* 2254GAT(689)* ; 2309GAT(706)
g676 and 2196GAT(656)* 2251GAT(690)* ; 2305GAT(707)
g677 and 2191GAT(659)* 2248GAT(691)* ; 2301GAT(708)
g678 and 2186GAT(662)* 2245GAT(692)* ; 2297GAT(709)
g679 and 2181GAT(665)* 2242GAT(693)* ; 2293GAT(710)
g680 and 2176GAT(668)* 2239GAT(694)* ; 2289GAT(711)
g681 and 2171GAT(671)* 2236GAT(695)* ; 2285GAT(712)
g682 and 2166GAT(674)* 2233GAT(696)* ; 2281GAT(713)
g683 and 2161GAT(677)* 2230GAT(697)* ; 2277GAT(714)
g684 and 2156GAT(680)* 2227GAT(698)* ; 2273GAT(715)
g685 and 2151GAT(682)* 2224GAT(699)* ; 2269GAT(716)
g686 and 2322GAT(703)* 2145GAT(623)* ; 2359GAT(717)
g687 and 2322GAT(703)* 2266GAT(684)* ; 2357GAT(718)
g688 and 2318GAT(704)* 2317GAT(702)* ; 2350GAT(719)
g689 and 2313GAT(705)* 2257GAT(688)* ; 2348GAT(720)
g690 and 1227GAT(59)* 2322GAT(703)* ; 2358GAT(721)
g691 and 2309GAT(706)* 2254GAT(689)* ; 2346GAT(722)
g692 and 1179GAT(75)* 2319GAT(701)* ; 2353GAT(723)
g693 and 2305GAT(707)* 2251GAT(690)* ; 2344GAT(724)
g694 and 2206GAT(650)* 2313GAT(705)* ; 2349GAT(725)
g695 and 2301GAT(708)* 2248GAT(691)* ; 2342GAT(726)
g696 and 2201GAT(653)* 2309GAT(706)* ; 2347GAT(727)
g697 and 2297GAT(709)* 2245GAT(692)* ; 2340GAT(728)
g698 and 2196GAT(656)* 2305GAT(707)* ; 2345GAT(729)
g699 and 2293GAT(710)* 2242GAT(693)* ; 2338GAT(730)
g700 and 2191GAT(659)* 2301GAT(708)* ; 2343GAT(731)
g701 and 2289GAT(711)* 2239GAT(694)* ; 2336GAT(732)
g702 and 2186GAT(662)* 2297GAT(709)* ; 2341GAT(733)
g703 and 2285GAT(712)* 2236GAT(695)* ; 2334GAT(734)
g704 and 2181GAT(665)* 2293GAT(710)* ; 2339GAT(735)
g705 and 2281GAT(713)* 2233GAT(696)* ; 2332GAT(736)
g706 and 2176GAT(668)* 2289GAT(711)* ; 2337GAT(737)
g707 and 2277GAT(714)* 2230GAT(697)* ; 2330GAT(738)
g708 and 2171GAT(671)* 2285GAT(712)* ; 2335GAT(739)
g709 and 2273GAT(715)* 2227GAT(698)* ; 2328GAT(740)
g710 and 2166GAT(674)* 2281GAT(713)* ; 2333GAT(741)
g711 and 2269GAT(716)* 2224GAT(699)* ; 2326GAT(742)
g712 and 2161GAT(677)* 2277GAT(714)* ; 2331GAT(743)
g713 and 2156GAT(680)* 2273GAT(715)* ; 2329GAT(744)
g714 and 2151GAT(682)* 2269GAT(716)* ; 2327GAT(745)
g715 and 2359GAT(717)* 1275GAT(43)* ; 2410GAT(746)
g716 and 2358GAT(721)* 2357GAT(718)* ; 2407GAT(747)
g717 and 2353GAT(723)* 2217GAT(643)* ; 2404GAT(748)
g718 and 2353GAT(723)* 2319GAT(701)* ; 2402GAT(749)
g719 and 2349GAT(725)* 2348GAT(720)* ; 2395GAT(750)
g720 and 2347GAT(727)* 2346GAT(722)* ; 2392GAT(751)
g721 and 1179GAT(75)* 2353GAT(723)* ; 2403GAT(752)
g722 and 2345GAT(729)* 2344GAT(724)* ; 2389GAT(753)
g723 and 1131GAT(91)* 2350GAT(719)* ; 2398GAT(754)
g724 and 2343GAT(731)* 2342GAT(726)* ; 2386GAT(755)
g725 and 2341GAT(733)* 2340GAT(728)* ; 2383GAT(756)
g726 and 2339GAT(735)* 2338GAT(730)* ; 2380GAT(757)
g727 and 2337GAT(737)* 2336GAT(732)* ; 2377GAT(758)
g728 and 2335GAT(739)* 2334GAT(734)* ; 2374GAT(759)
g729 and 2333GAT(741)* 2332GAT(736)* ; 2371GAT(760)
g730 and 2331GAT(743)* 2330GAT(738)* ; 2368GAT(761)
g731 and 2329GAT(744)* 2328GAT(740)* ; 2365GAT(762)
g732 and 2327GAT(745)* 2326GAT(742)* ; 2362GAT(763)
g733 and 2410GAT(746)* 1275GAT(43)* ; 2474GAT(764)
g734 and 2359GAT(717)* 2410GAT(746)* ; 2475GAT(765)
g735 and 2404GAT(748)* 2407GAT(747)* ; 2470GAT(766)
g736 and 2403GAT(752)* 2402GAT(749)* ; 2467GAT(767)
g737 and 2398GAT(754)* 2260GAT(687)* ; 2464GAT(768)
g738 and 2398GAT(754)* 2350GAT(719)* ; 2462GAT(769)
g739 and 1131GAT(91)* 2398GAT(754)* ; 2463GAT(770)
g740 and 1083GAT(107)* 2395GAT(750)* ; 2458GAT(771)
g741 and 1035GAT(123)* 2392GAT(751)* ; 2454GAT(772)
g742 and 987GAT(139)* 2389GAT(753)* ; 2450GAT(773)
g743 and 939GAT(155)* 2386GAT(755)* ; 2446GAT(774)
g744 and 891GAT(171)* 2383GAT(756)* ; 2442GAT(775)
g745 and 843GAT(187)* 2380GAT(757)* ; 2438GAT(776)
g746 and 795GAT(203)* 2377GAT(758)* ; 2434GAT(777)
g747 and 747GAT(219)* 2374GAT(759)* ; 2430GAT(778)
g748 and 699GAT(235)* 2371GAT(760)* ; 2426GAT(779)
g749 and 651GAT(251)* 2368GAT(761)* ; 2422GAT(780)
g750 and 603GAT(267)* 2365GAT(762)* ; 2418GAT(781)
g751 and 555GAT(283)* 2362GAT(763)* ; 2414GAT(782)
g752 and 2475GAT(765)* 2474GAT(764)* ; 2545GAT(783)
g753 and 2470GAT(766)* 2407GAT(747)* ; 2543GAT(784)
g754 and 2404GAT(748)* 2470GAT(766)* ; 2544GAT(785)
g755 and 2464GAT(768)* 2467GAT(767)* ; 2539GAT(786)
g756 and 2463GAT(770)* 2462GAT(769)* ; 2536GAT(787)
g757 and 2458GAT(771)* 2395GAT(750)* ; 2531GAT(788)
g758 and 2454GAT(772)* 2392GAT(751)* ; 2526GAT(789)
g759 and 2450GAT(773)* 2389GAT(753)* ; 2521GAT(790)
g760 and 2458GAT(771)* 2313GAT(705)* ; 2533GAT(791)
g761 and 2446GAT(774)* 2386GAT(755)* ; 2516GAT(792)
g762 and 1083GAT(107)* 2458GAT(771)* ; 2532GAT(793)
g763 and 2454GAT(772)* 2309GAT(706)* ; 2528GAT(794)
g764 and 2442GAT(775)* 2383GAT(756)* ; 2511GAT(795)
g765 and 1035GAT(123)* 2454GAT(772)* ; 2527GAT(796)
g766 and 2450GAT(773)* 2305GAT(707)* ; 2523GAT(797)
g767 and 2438GAT(776)* 2380GAT(757)* ; 2506GAT(798)
g768 and 987GAT(139)* 2450GAT(773)* ; 2522GAT(799)
g769 and 2446GAT(774)* 2301GAT(708)* ; 2518GAT(800)
g770 and 2434GAT(777)* 2377GAT(758)* ; 2501GAT(801)
g771 and 939GAT(155)* 2446GAT(774)* ; 2517GAT(802)
g772 and 2442GAT(775)* 2297GAT(709)* ; 2513GAT(803)
g773 and 2430GAT(778)* 2374GAT(759)* ; 2496GAT(804)
g774 and 891GAT(171)* 2442GAT(775)* ; 2512GAT(805)
g775 and 2438GAT(776)* 2293GAT(710)* ; 2508GAT(806)
g776 and 2426GAT(779)* 2371GAT(760)* ; 2491GAT(807)
g777 and 843GAT(187)* 2438GAT(776)* ; 2507GAT(808)
g778 and 2434GAT(777)* 2289GAT(711)* ; 2503GAT(809)
g779 and 2422GAT(780)* 2368GAT(761)* ; 2486GAT(810)
g780 and 795GAT(203)* 2434GAT(777)* ; 2502GAT(811)
g781 and 2430GAT(778)* 2285GAT(712)* ; 2498GAT(812)
g782 and 2418GAT(781)* 2365GAT(762)* ; 2481GAT(813)
g783 and 747GAT(219)* 2430GAT(778)* ; 2497GAT(814)
g784 and 2426GAT(779)* 2281GAT(713)* ; 2493GAT(815)
g785 and 2414GAT(782)* 2362GAT(763)* ; 2476GAT(816)
g786 and 699GAT(235)* 2426GAT(779)* ; 2492GAT(817)
g787 and 2422GAT(780)* 2277GAT(714)* ; 2488GAT(818)
g788 and 651GAT(251)* 2422GAT(780)* ; 2487GAT(819)
g789 and 2418GAT(781)* 2273GAT(715)* ; 2483GAT(820)
g790 and 603GAT(267)* 2418GAT(781)* ; 2482GAT(821)
g791 and 2414GAT(782)* 2269GAT(716)* ; 2478GAT(822)
g792 and 555GAT(283)* 2414GAT(782)* ; 2477GAT(823)
g793 and 2544GAT(785)* 2543GAT(784)* ; 2588GAT(824)
g794 and 2539GAT(786)* 2467GAT(767)* ; 2586GAT(825)
g795 and 2464GAT(768)* 2539GAT(786)* ; 2587GAT(826)
g796 and 2533GAT(791)* 2536GAT(787)* ; 2582GAT(827)
g797 and 2532GAT(793)* 2531GAT(788)* ; 2579GAT(828)
g798 and 1230GAT(58)* 2545GAT(783)* ; 2591GAT(829)
g799 and 2527GAT(796)* 2526GAT(789)* ; 2576GAT(830)
g800 and 2522GAT(799)* 2521GAT(790)* ; 2573GAT(831)
g801 and 2517GAT(802)* 2516GAT(792)* ; 2570GAT(832)
g802 and 2512GAT(805)* 2511GAT(795)* ; 2567GAT(833)
g803 and 2507GAT(808)* 2506GAT(798)* ; 2564GAT(834)
g804 and 2502GAT(811)* 2501GAT(801)* ; 2561GAT(835)
g805 and 2497GAT(814)* 2496GAT(804)* ; 2558GAT(836)
g806 and 2492GAT(817)* 2491GAT(807)* ; 2555GAT(837)
g807 and 2487GAT(819)* 2486GAT(810)* ; 2552GAT(838)
g808 and 2482GAT(821)* 2481GAT(813)* ; 2549GAT(839)
g809 and 2477GAT(823)* 2476GAT(816)* ; 2548GAT(840)
g810 and 2591GAT(829)* 2410GAT(746)* ; 2650GAT(841)
g811 and 2591GAT(829)* 2545GAT(783)* ; 2648GAT(842)
g812 and 2587GAT(826)* 2586GAT(825)* ; 2641GAT(843)
g813 and 2582GAT(827)* 2536GAT(787)* ; 2639GAT(844)
g814 and 1230GAT(58)* 2591GAT(829)* ; 2649GAT(845)
g815 and 1182GAT(74)* 2588GAT(824)* ; 2644GAT(846)
g816 and 2533GAT(791)* 2582GAT(827)* ; 2640GAT(847)
g817 and 2528GAT(794)* 2579GAT(828)* ; 2635GAT(848)
g818 and 2523GAT(797)* 2576GAT(830)* ; 2631GAT(849)
g819 and 2518GAT(800)* 2573GAT(831)* ; 2627GAT(850)
g820 and 2513GAT(803)* 2570GAT(832)* ; 2623GAT(851)
g821 and 2508GAT(806)* 2567GAT(833)* ; 2619GAT(852)
g822 and 2503GAT(809)* 2564GAT(834)* ; 2615GAT(853)
g823 and 2498GAT(812)* 2561GAT(835)* ; 2611GAT(854)
g824 and 2493GAT(815)* 2558GAT(836)* ; 2607GAT(855)
g825 and 2488GAT(818)* 2555GAT(837)* ; 2603GAT(856)
g826 and 2483GAT(820)* 2552GAT(838)* ; 2599GAT(857)
g827 and 2478GAT(822)* 2549GAT(839)* ; 2595GAT(858)
g828 and 2650GAT(841)* 1278GAT(42)* ; 2690GAT(859)
g829 and 2649GAT(845)* 2648GAT(842)* ; 2687GAT(860)
g830 and 2644GAT(846)* 2470GAT(766)* ; 2684GAT(861)
g831 and 2644GAT(846)* 2588GAT(824)* ; 2682GAT(862)
g832 and 2640GAT(847)* 2639GAT(844)* ; 2675GAT(863)
g833 and 2635GAT(848)* 2579GAT(828)* ; 2673GAT(864)
g834 and 2631GAT(849)* 2576GAT(830)* ; 2671GAT(865)
g835 and 1182GAT(74)* 2644GAT(846)* ; 2683GAT(866)
g836 and 2627GAT(850)* 2573GAT(831)* ; 2669GAT(867)
g837 and 1134GAT(90)* 2641GAT(843)* ; 2678GAT(868)
g838 and 2623GAT(851)* 2570GAT(832)* ; 2667GAT(869)
g839 and 2528GAT(794)* 2635GAT(848)* ; 2674GAT(870)
g840 and 2619GAT(852)* 2567GAT(833)* ; 2665GAT(871)
g841 and 2523GAT(797)* 2631GAT(849)* ; 2672GAT(872)
g842 and 2615GAT(853)* 2564GAT(834)* ; 2663GAT(873)
g843 and 2518GAT(800)* 2627GAT(850)* ; 2670GAT(874)
g844 and 2611GAT(854)* 2561GAT(835)* ; 2661GAT(875)
g845 and 2513GAT(803)* 2623GAT(851)* ; 2668GAT(876)
g846 and 2607GAT(855)* 2558GAT(836)* ; 2659GAT(877)
g847 and 2508GAT(806)* 2619GAT(852)* ; 2666GAT(878)
g848 and 2603GAT(856)* 2555GAT(837)* ; 2657GAT(879)
g849 and 2503GAT(809)* 2615GAT(853)* ; 2664GAT(880)
g850 and 2599GAT(857)* 2552GAT(838)* ; 2655GAT(881)
g851 and 2498GAT(812)* 2611GAT(854)* ; 2662GAT(882)
g852 and 2595GAT(858)* 2549GAT(839)* ; 2653GAT(883)
g853 and 2493GAT(815)* 2607GAT(855)* ; 2660GAT(884)
g854 and 2488GAT(818)* 2603GAT(856)* ; 2658GAT(885)
g855 and 2483GAT(820)* 2599GAT(857)* ; 2656GAT(886)
g856 and 2478GAT(822)* 2595GAT(858)* ; 2654GAT(887)
g857 and 2690GAT(859)* 1278GAT(42)* ; 2743GAT(888)
g858 and 2650GAT(841)* 2690GAT(859)* ; 2744GAT(889)
g859 and 2684GAT(861)* 2687GAT(860)* ; 2739GAT(890)
g860 and 2683GAT(866)* 2682GAT(862)* ; 2736GAT(891)
g861 and 2678GAT(868)* 2539GAT(786)* ; 2733GAT(892)
g862 and 2678GAT(868)* 2641GAT(843)* ; 2731GAT(893)
g863 and 2674GAT(870)* 2673GAT(864)* ; 2724GAT(894)
g864 and 2672GAT(872)* 2671GAT(865)* ; 2721GAT(895)
g865 and 2670GAT(874)* 2669GAT(867)* ; 2718GAT(896)
g866 and 1134GAT(90)* 2678GAT(868)* ; 2732GAT(897)
g867 and 2668GAT(876)* 2667GAT(869)* ; 2715GAT(898)
g868 and 1086GAT(106)* 2675GAT(863)* ; 2727GAT(899)
g869 and 2666GAT(878)* 2665GAT(871)* ; 2712GAT(900)
g870 and 2664GAT(880)* 2663GAT(873)* ; 2709GAT(901)
g871 and 2662GAT(882)* 2661GAT(875)* ; 2706GAT(902)
g872 and 2660GAT(884)* 2659GAT(877)* ; 2703GAT(903)
g873 and 2658GAT(885)* 2657GAT(879)* ; 2700GAT(904)
g874 and 2656GAT(886)* 2655GAT(881)* ; 2697GAT(905)
g875 and 2654GAT(887)* 2653GAT(883)* ; 2694GAT(906)
g876 and 2744GAT(889)* 2743GAT(888)* ; 2803GAT(907)
g877 and 2739GAT(890)* 2687GAT(860)* ; 2801GAT(908)
g878 and 2684GAT(861)* 2739GAT(890)* ; 2802GAT(909)
g879 and 2733GAT(892)* 2736GAT(891)* ; 2797GAT(910)
g880 and 2732GAT(897)* 2731GAT(893)* ; 2794GAT(911)
g881 and 2727GAT(899)* 2582GAT(827)* ; 2791GAT(912)
g882 and 2727GAT(899)* 2675GAT(863)* ; 2789GAT(913)
g883 and 1086GAT(106)* 2727GAT(899)* ; 2790GAT(914)
g884 and 1038GAT(122)* 2724GAT(894)* ; 2785GAT(915)
g885 and 990GAT(138)* 2721GAT(895)* ; 2781GAT(916)
g886 and 942GAT(154)* 2718GAT(896)* ; 2777GAT(917)
g887 and 894GAT(170)* 2715GAT(898)* ; 2773GAT(918)
g888 and 846GAT(186)* 2712GAT(900)* ; 2769GAT(919)
g889 and 798GAT(202)* 2709GAT(901)* ; 2765GAT(920)
g890 and 750GAT(218)* 2706GAT(902)* ; 2761GAT(921)
g891 and 702GAT(234)* 2703GAT(903)* ; 2757GAT(922)
g892 and 654GAT(250)* 2700GAT(904)* ; 2753GAT(923)
g893 and 606GAT(266)* 2697GAT(905)* ; 2749GAT(924)
g894 and 558GAT(282)* 2694GAT(906)* ; 2745GAT(925)
g895 and 2802GAT(909)* 2801GAT(908)* ; 2870GAT(926)
g896 and 2797GAT(910)* 2736GAT(891)* ; 2868GAT(927)
g897 and 2733GAT(892)* 2797GAT(910)* ; 2869GAT(928)
g898 and 2791GAT(912)* 2794GAT(911)* ; 2864GAT(929)
g899 and 2790GAT(914)* 2789GAT(913)* ; 2861GAT(930)
g900 and 2785GAT(915)* 2724GAT(894)* ; 2856GAT(931)
g901 and 1233GAT(57)* 2803GAT(907)* ; 2873GAT(932)
g902 and 2781GAT(916)* 2721GAT(895)* ; 2851GAT(933)
g903 and 2777GAT(917)* 2718GAT(896)* ; 2846GAT(934)
g904 and 2773GAT(918)* 2715GAT(898)* ; 2841GAT(935)
g905 and 2785GAT(915)* 2635GAT(848)* ; 2858GAT(936)
g906 and 2769GAT(919)* 2712GAT(900)* ; 2836GAT(937)
g907 and 1038GAT(122)* 2785GAT(915)* ; 2857GAT(938)
g908 and 2781GAT(916)* 2631GAT(849)* ; 2853GAT(939)
g909 and 2765GAT(920)* 2709GAT(901)* ; 2831GAT(940)
g910 and 990GAT(138)* 2781GAT(916)* ; 2852GAT(941)
g911 and 2777GAT(917)* 2627GAT(850)* ; 2848GAT(942)
g912 and 2761GAT(921)* 2706GAT(902)* ; 2826GAT(943)
g913 and 942GAT(154)* 2777GAT(917)* ; 2847GAT(944)
g914 and 2773GAT(918)* 2623GAT(851)* ; 2843GAT(945)
g915 and 2757GAT(922)* 2703GAT(903)* ; 2821GAT(946)
g916 and 894GAT(170)* 2773GAT(918)* ; 2842GAT(947)
g917 and 2769GAT(919)* 2619GAT(852)* ; 2838GAT(948)
g918 and 2753GAT(923)* 2700GAT(904)* ; 2816GAT(949)
g919 and 846GAT(186)* 2769GAT(919)* ; 2837GAT(950)
g920 and 2765GAT(920)* 2615GAT(853)* ; 2833GAT(951)
g921 and 2749GAT(924)* 2697GAT(905)* ; 2811GAT(952)
g922 and 798GAT(202)* 2765GAT(920)* ; 2832GAT(953)
g923 and 2761GAT(921)* 2611GAT(854)* ; 2828GAT(954)
g924 and 2745GAT(925)* 2694GAT(906)* ; 2806GAT(955)
g925 and 750GAT(218)* 2761GAT(921)* ; 2827GAT(956)
g926 and 2757GAT(922)* 2607GAT(855)* ; 2823GAT(957)
g927 and 702GAT(234)* 2757GAT(922)* ; 2822GAT(958)
g928 and 2753GAT(923)* 2603GAT(856)* ; 2818GAT(959)
g929 and 654GAT(250)* 2753GAT(923)* ; 2817GAT(960)
g930 and 2749GAT(924)* 2599GAT(857)* ; 2813GAT(961)
g931 and 606GAT(266)* 2749GAT(924)* ; 2812GAT(962)
g932 and 2745GAT(925)* 2595GAT(858)* ; 2808GAT(963)
g933 and 558GAT(282)* 2745GAT(925)* ; 2807GAT(964)
g934 and 2873GAT(932)* 2690GAT(859)* ; 2923GAT(965)
g935 and 2873GAT(932)* 2803GAT(907)* ; 2921GAT(966)
g936 and 2869GAT(928)* 2868GAT(927)* ; 2914GAT(967)
g937 and 2864GAT(929)* 2794GAT(911)* ; 2912GAT(968)
g938 and 2791GAT(912)* 2864GAT(929)* ; 2913GAT(969)
g939 and 2858GAT(936)* 2861GAT(930)* ; 2908GAT(970)
g940 and 2857GAT(938)* 2856GAT(931)* ; 2905GAT(971)
g941 and 1233GAT(57)* 2873GAT(932)* ; 2922GAT(972)
g942 and 2852GAT(941)* 2851GAT(933)* ; 2902GAT(973)
g943 and 1185GAT(73)* 2870GAT(926)* ; 2917GAT(974)
g944 and 2847GAT(944)* 2846GAT(934)* ; 2899GAT(975)
g945 and 2842GAT(947)* 2841GAT(935)* ; 2896GAT(976)
g946 and 2837GAT(950)* 2836GAT(937)* ; 2893GAT(977)
g947 and 2832GAT(953)* 2831GAT(940)* ; 2890GAT(978)
g948 and 2827GAT(956)* 2826GAT(943)* ; 2887GAT(979)
g949 and 2822GAT(958)* 2821GAT(946)* ; 2884GAT(980)
g950 and 2817GAT(960)* 2816GAT(949)* ; 2881GAT(981)
g951 and 2812GAT(962)* 2811GAT(952)* ; 2878GAT(982)
g952 and 2807GAT(964)* 2806GAT(955)* ; 2877GAT(983)
g953 and 2923GAT(965)* 1281GAT(41)* ; 2983GAT(984)
g954 and 2922GAT(972)* 2921GAT(966)* ; 2980GAT(985)
g955 and 2917GAT(974)* 2739GAT(890)* ; 2977GAT(986)
g956 and 2917GAT(974)* 2870GAT(926)* ; 2975GAT(987)
g957 and 2913GAT(969)* 2912GAT(968)* ; 2968GAT(988)
g958 and 2908GAT(970)* 2861GAT(930)* ; 2966GAT(989)
g959 and 1185GAT(73)* 2917GAT(974)* ; 2976GAT(990)
g960 and 1137GAT(89)* 2914GAT(967)* ; 2971GAT(991)
g961 and 2858GAT(936)* 2908GAT(970)* ; 2967GAT(992)
g962 and 2853GAT(939)* 2905GAT(971)* ; 2962GAT(993)
g963 and 2848GAT(942)* 2902GAT(973)* ; 2958GAT(994)
g964 and 2843GAT(945)* 2899GAT(975)* ; 2954GAT(995)
g965 and 2838GAT(948)* 2896GAT(976)* ; 2950GAT(996)
g966 and 2833GAT(951)* 2893GAT(977)* ; 2946GAT(997)
g967 and 2828GAT(954)* 2890GAT(978)* ; 2942GAT(998)
g968 and 2823GAT(957)* 2887GAT(979)* ; 2938GAT(999)
g969 and 2818GAT(959)* 2884GAT(980)* ; 2934GAT(1000)
g970 and 2813GAT(961)* 2881GAT(981)* ; 2930GAT(1001)
g971 and 2808GAT(963)* 2878GAT(982)* ; 2926GAT(1002)
g972 and 2983GAT(984)* 1281GAT(41)* ; 3026GAT(1003)
g973 and 2923GAT(965)* 2983GAT(984)* ; 3027GAT(1004)
g974 and 2977GAT(986)* 2980GAT(985)* ; 3022GAT(1005)
g975 and 2976GAT(990)* 2975GAT(987)* ; 3019GAT(1006)
g976 and 2971GAT(991)* 2797GAT(910)* ; 3016GAT(1007)
g977 and 2971GAT(991)* 2914GAT(967)* ; 3014GAT(1008)
g978 and 2967GAT(992)* 2966GAT(989)* ; 3007GAT(1009)
g979 and 2962GAT(993)* 2905GAT(971)* ; 3005GAT(1010)
g980 and 2958GAT(994)* 2902GAT(973)* ; 3003GAT(1011)
g981 and 2954GAT(995)* 2899GAT(975)* ; 3001GAT(1012)
g982 and 1137GAT(89)* 2971GAT(991)* ; 3015GAT(1013)
g983 and 2950GAT(996)* 2896GAT(976)* ; 2999GAT(1014)
g984 and 1089GAT(105)* 2968GAT(988)* ; 3010GAT(1015)
g985 and 2946GAT(997)* 2893GAT(977)* ; 2997GAT(1016)
g986 and 2853GAT(939)* 2962GAT(993)* ; 3006GAT(1017)
g987 and 2942GAT(998)* 2890GAT(978)* ; 2995GAT(1018)
g988 and 2848GAT(942)* 2958GAT(994)* ; 3004GAT(1019)
g989 and 2938GAT(999)* 2887GAT(979)* ; 2993GAT(1020)
g990 and 2843GAT(945)* 2954GAT(995)* ; 3002GAT(1021)
g991 and 2934GAT(1000)* 2884GAT(980)* ; 2991GAT(1022)
g992 and 2838GAT(948)* 2950GAT(996)* ; 3000GAT(1023)
g993 and 2930GAT(1001)* 2881GAT(981)* ; 2989GAT(1024)
g994 and 2833GAT(951)* 2946GAT(997)* ; 2998GAT(1025)
g995 and 2926GAT(1002)* 2878GAT(982)* ; 2987GAT(1026)
g996 and 2828GAT(954)* 2942GAT(998)* ; 2996GAT(1027)
g997 and 2823GAT(957)* 2938GAT(999)* ; 2994GAT(1028)
g998 and 2818GAT(959)* 2934GAT(1000)* ; 2992GAT(1029)
g999 and 2813GAT(961)* 2930GAT(1001)* ; 2990GAT(1030)
g1000 and 2808GAT(963)* 2926GAT(1002)* ; 2988GAT(1031)
g1001 and 3027GAT(1004)* 3026GAT(1003)* ; 3076GAT(1032)
g1002 and 3022GAT(1005)* 2980GAT(985)* ; 3074GAT(1033)
g1003 and 2977GAT(986)* 3022GAT(1005)* ; 3075GAT(1034)
g1004 and 3016GAT(1007)* 3019GAT(1006)* ; 3070GAT(1035)
g1005 and 3015GAT(1013)* 3014GAT(1008)* ; 3067GAT(1036)
g1006 and 3010GAT(1015)* 2864GAT(929)* ; 3064GAT(1037)
g1007 and 3010GAT(1015)* 2968GAT(988)* ; 3062GAT(1038)
g1008 and 3006GAT(1017)* 3005GAT(1010)* ; 3055GAT(1039)
g1009 and 3004GAT(1019)* 3003GAT(1011)* ; 3052GAT(1040)
g1010 and 3002GAT(1021)* 3001GAT(1012)* ; 3049GAT(1041)
g1011 and 3000GAT(1023)* 2999GAT(1014)* ; 3046GAT(1042)
g1012 and 1089GAT(105)* 3010GAT(1015)* ; 3063GAT(1043)
g1013 and 2998GAT(1025)* 2997GAT(1016)* ; 3043GAT(1044)
g1014 and 1041GAT(121)* 3007GAT(1009)* ; 3058GAT(1045)
g1015 and 2996GAT(1027)* 2995GAT(1018)* ; 3040GAT(1046)
g1016 and 2994GAT(1028)* 2993GAT(1020)* ; 3037GAT(1047)
g1017 and 2992GAT(1029)* 2991GAT(1022)* ; 3034GAT(1048)
g1018 and 2990GAT(1030)* 2989GAT(1024)* ; 3031GAT(1049)
g1019 and 2988GAT(1031)* 2987GAT(1026)* ; 3028GAT(1050)
g1020 and 3075GAT(1034)* 3074GAT(1033)* ; 3133GAT(1051)
g1021 and 3070GAT(1035)* 3019GAT(1006)* ; 3131GAT(1052)
g1022 and 3016GAT(1007)* 3070GAT(1035)* ; 3132GAT(1053)
g1023 and 3064GAT(1037)* 3067GAT(1036)* ; 3127GAT(1054)
g1024 and 3063GAT(1043)* 3062GAT(1038)* ; 3124GAT(1055)
g1025 and 3058GAT(1045)* 2908GAT(970)* ; 3121GAT(1056)
g1026 and 3058GAT(1045)* 3007GAT(1009)* ; 3119GAT(1057)
g1027 and 1236GAT(56)* 3076GAT(1032)* ; 3136GAT(1058)
g1028 and 1041GAT(121)* 3058GAT(1045)* ; 3120GAT(1059)
g1029 and 993GAT(137)* 3055GAT(1039)* ; 3115GAT(1060)
g1030 and 945GAT(153)* 3052GAT(1040)* ; 3111GAT(1061)
g1031 and 897GAT(169)* 3049GAT(1041)* ; 3107GAT(1062)
g1032 and 849GAT(185)* 3046GAT(1042)* ; 3103GAT(1063)
g1033 and 801GAT(201)* 3043GAT(1044)* ; 3099GAT(1064)
g1034 and 753GAT(217)* 3040GAT(1046)* ; 3095GAT(1065)
g1035 and 705GAT(233)* 3037GAT(1047)* ; 3091GAT(1066)
g1036 and 657GAT(249)* 3034GAT(1048)* ; 3087GAT(1067)
g1037 and 609GAT(265)* 3031GAT(1049)* ; 3083GAT(1068)
g1038 and 561GAT(281)* 3028GAT(1050)* ; 3079GAT(1069)
g1039 and 3136GAT(1058)* 2983GAT(984)* ; 3208GAT(1070)
g1040 and 3136GAT(1058)* 3076GAT(1032)* ; 3206GAT(1071)
g1041 and 3132GAT(1053)* 3131GAT(1052)* ; 3199GAT(1072)
g1042 and 3127GAT(1054)* 3067GAT(1036)* ; 3197GAT(1073)
g1043 and 3064GAT(1037)* 3127GAT(1054)* ; 3198GAT(1074)
g1044 and 3121GAT(1056)* 3124GAT(1055)* ; 3193GAT(1075)
g1045 and 3120GAT(1059)* 3119GAT(1057)* ; 3190GAT(1076)
g1046 and 3115GAT(1060)* 3055GAT(1039)* ; 3185GAT(1077)
g1047 and 1236GAT(56)* 3136GAT(1058)* ; 3207GAT(1078)
g1048 and 3111GAT(1061)* 3052GAT(1040)* ; 3180GAT(1079)
g1049 and 1188GAT(72)* 3133GAT(1051)* ; 3202GAT(1080)
g1050 and 3107GAT(1062)* 3049GAT(1041)* ; 3175GAT(1081)
g1051 and 3103GAT(1063)* 3046GAT(1042)* ; 3170GAT(1082)
g1052 and 3099GAT(1064)* 3043GAT(1044)* ; 3165GAT(1083)
g1053 and 3115GAT(1060)* 2962GAT(993)* ; 3187GAT(1084)
g1054 and 3095GAT(1065)* 3040GAT(1046)* ; 3160GAT(1085)
g1055 and 993GAT(137)* 3115GAT(1060)* ; 3186GAT(1086)
g1056 and 3111GAT(1061)* 2958GAT(994)* ; 3182GAT(1087)
g1057 and 3091GAT(1066)* 3037GAT(1047)* ; 3155GAT(1088)
g1058 and 945GAT(153)* 3111GAT(1061)* ; 3181GAT(1089)
g1059 and 3107GAT(1062)* 2954GAT(995)* ; 3177GAT(1090)
g1060 and 3087GAT(1067)* 3034GAT(1048)* ; 3150GAT(1091)
g1061 and 897GAT(169)* 3107GAT(1062)* ; 3176GAT(1092)
g1062 and 3103GAT(1063)* 2950GAT(996)* ; 3172GAT(1093)
g1063 and 3083GAT(1068)* 3031GAT(1049)* ; 3145GAT(1094)
g1064 and 849GAT(185)* 3103GAT(1063)* ; 3171GAT(1095)
g1065 and 3099GAT(1064)* 2946GAT(997)* ; 3167GAT(1096)
g1066 and 3079GAT(1069)* 3028GAT(1050)* ; 3140GAT(1097)
g1067 and 801GAT(201)* 3099GAT(1064)* ; 3166GAT(1098)
g1068 and 3095GAT(1065)* 2942GAT(998)* ; 3162GAT(1099)
g1069 and 753GAT(217)* 3095GAT(1065)* ; 3161GAT(1100)
g1070 and 3091GAT(1066)* 2938GAT(999)* ; 3157GAT(1101)
g1071 and 705GAT(233)* 3091GAT(1066)* ; 3156GAT(1102)
g1072 and 3087GAT(1067)* 2934GAT(1000)* ; 3152GAT(1103)
g1073 and 657GAT(249)* 3087GAT(1067)* ; 3151GAT(1104)
g1074 and 3083GAT(1068)* 2930GAT(1001)* ; 3147GAT(1105)
g1075 and 609GAT(265)* 3083GAT(1068)* ; 3146GAT(1106)
g1076 and 3079GAT(1069)* 2926GAT(1002)* ; 3142GAT(1107)
g1077 and 561GAT(281)* 3079GAT(1069)* ; 3141GAT(1108)
g1078 and 3208GAT(1070)* 1284GAT(40)* ; 3260GAT(1109)
g1079 and 3207GAT(1078)* 3206GAT(1071)* ; 3257GAT(1110)
g1080 and 3202GAT(1080)* 3022GAT(1005)* ; 3254GAT(1111)
g1081 and 3202GAT(1080)* 3133GAT(1051)* ; 3252GAT(1112)
g1082 and 3198GAT(1074)* 3197GAT(1073)* ; 3245GAT(1113)
g1083 and 3193GAT(1075)* 3124GAT(1055)* ; 3243GAT(1114)
g1084 and 3121GAT(1056)* 3193GAT(1075)* ; 3244GAT(1115)
g1085 and 3187GAT(1084)* 3190GAT(1076)* ; 3239GAT(1116)
g1086 and 3186GAT(1086)* 3185GAT(1077)* ; 3236GAT(1117)
g1087 and 3181GAT(1089)* 3180GAT(1079)* ; 3233GAT(1118)
g1088 and 1188GAT(72)* 3202GAT(1080)* ; 3253GAT(1119)
g1089 and 3176GAT(1092)* 3175GAT(1081)* ; 3230GAT(1120)
g1090 and 1140GAT(88)* 3199GAT(1072)* ; 3248GAT(1121)
g1091 and 3171GAT(1095)* 3170GAT(1082)* ; 3227GAT(1122)
g1092 and 3166GAT(1098)* 3165GAT(1083)* ; 3224GAT(1123)
g1093 and 3161GAT(1100)* 3160GAT(1085)* ; 3221GAT(1124)
g1094 and 3156GAT(1102)* 3155GAT(1088)* ; 3218GAT(1125)
g1095 and 3151GAT(1104)* 3150GAT(1091)* ; 3215GAT(1126)
g1096 and 3146GAT(1106)* 3145GAT(1094)* ; 3212GAT(1127)
g1097 and 3141GAT(1108)* 3140GAT(1097)* ; 3211GAT(1128)
g1098 and 3260GAT(1109)* 1284GAT(40)* ; 3321GAT(1129)
g1099 and 3208GAT(1070)* 3260GAT(1109)* ; 3322GAT(1130)
g1100 and 3254GAT(1111)* 3257GAT(1110)* ; 3317GAT(1131)
g1101 and 3253GAT(1119)* 3252GAT(1112)* ; 3314GAT(1132)
g1102 and 3248GAT(1121)* 3070GAT(1035)* ; 3311GAT(1133)
g1103 and 3248GAT(1121)* 3199GAT(1072)* ; 3309GAT(1134)
g1104 and 3244GAT(1115)* 3243GAT(1114)* ; 3302GAT(1135)
g1105 and 3239GAT(1116)* 3190GAT(1076)* ; 3300GAT(1136)
g1106 and 1140GAT(88)* 3248GAT(1121)* ; 3310GAT(1137)
g1107 and 1092GAT(104)* 3245GAT(1113)* ; 3305GAT(1138)
g1108 and 3187GAT(1084)* 3239GAT(1116)* ; 3301GAT(1139)
g1109 and 3182GAT(1087)* 3236GAT(1117)* ; 3296GAT(1140)
g1110 and 3177GAT(1090)* 3233GAT(1118)* ; 3292GAT(1141)
g1111 and 3172GAT(1093)* 3230GAT(1120)* ; 3288GAT(1142)
g1112 and 3167GAT(1096)* 3227GAT(1122)* ; 3284GAT(1143)
g1113 and 3162GAT(1099)* 3224GAT(1123)* ; 3280GAT(1144)
g1114 and 3157GAT(1101)* 3221GAT(1124)* ; 3276GAT(1145)
g1115 and 3152GAT(1103)* 3218GAT(1125)* ; 3272GAT(1146)
g1116 and 3147GAT(1105)* 3215GAT(1126)* ; 3268GAT(1147)
g1117 and 3142GAT(1107)* 3212GAT(1127)* ; 3264GAT(1148)
g1118 and 3322GAT(1130)* 3321GAT(1129)* ; 3362GAT(1149)
g1119 and 3317GAT(1131)* 3257GAT(1110)* ; 3360GAT(1150)
g1120 and 3254GAT(1111)* 3317GAT(1131)* ; 3361GAT(1151)
g1121 and 3311GAT(1133)* 3314GAT(1132)* ; 3356GAT(1152)
g1122 and 3310GAT(1137)* 3309GAT(1134)* ; 3353GAT(1153)
g1123 and 3305GAT(1138)* 3127GAT(1054)* ; 3350GAT(1154)
g1124 and 3305GAT(1138)* 3245GAT(1113)* ; 3348GAT(1155)
g1125 and 3301GAT(1139)* 3300GAT(1136)* ; 3341GAT(1156)
g1126 and 3296GAT(1140)* 3236GAT(1117)* ; 3339GAT(1157)
g1127 and 3292GAT(1141)* 3233GAT(1118)* ; 3337GAT(1158)
g1128 and 3288GAT(1142)* 3230GAT(1120)* ; 3335GAT(1159)
g1129 and 3284GAT(1143)* 3227GAT(1122)* ; 3333GAT(1160)
g1130 and 1092GAT(104)* 3305GAT(1138)* ; 3349GAT(1161)
g1131 and 3280GAT(1144)* 3224GAT(1123)* ; 3331GAT(1162)
g1132 and 1044GAT(120)* 3302GAT(1135)* ; 3344GAT(1163)
g1133 and 3276GAT(1145)* 3221GAT(1124)* ; 3329GAT(1164)
g1134 and 3182GAT(1087)* 3296GAT(1140)* ; 3340GAT(1165)
g1135 and 3272GAT(1146)* 3218GAT(1125)* ; 3327GAT(1166)
g1136 and 3177GAT(1090)* 3292GAT(1141)* ; 3338GAT(1167)
g1137 and 3268GAT(1147)* 3215GAT(1126)* ; 3325GAT(1168)
g1138 and 3172GAT(1093)* 3288GAT(1142)* ; 3336GAT(1169)
g1139 and 3264GAT(1148)* 3212GAT(1127)* ; 3323GAT(1170)
g1140 and 3167GAT(1096)* 3284GAT(1143)* ; 3334GAT(1171)
g1141 and 3162GAT(1099)* 3280GAT(1144)* ; 3332GAT(1172)
g1142 and 3157GAT(1101)* 3276GAT(1145)* ; 3330GAT(1173)
g1143 and 3152GAT(1103)* 3272GAT(1146)* ; 3328GAT(1174)
g1144 and 3147GAT(1105)* 3268GAT(1147)* ; 3326GAT(1175)
g1145 and 3142GAT(1107)* 3264GAT(1148)* ; 3324GAT(1176)
g1146 and 3361GAT(1151)* 3360GAT(1150)* ; 3410GAT(1177)
g1147 and 3356GAT(1152)* 3314GAT(1132)* ; 3408GAT(1178)
g1148 and 3311GAT(1133)* 3356GAT(1152)* ; 3409GAT(1179)
g1149 and 3350GAT(1154)* 3353GAT(1153)* ; 3404GAT(1180)
g1150 and 3349GAT(1161)* 3348GAT(1155)* ; 3401GAT(1181)
g1151 and 3344GAT(1163)* 3193GAT(1075)* ; 3398GAT(1182)
g1152 and 3344GAT(1163)* 3302GAT(1135)* ; 3396GAT(1183)
g1153 and 3340GAT(1165)* 3339GAT(1157)* ; 3389GAT(1184)
g1154 and 1239GAT(55)* 3362GAT(1149)* ; 3413GAT(1185)
g1155 and 3338GAT(1167)* 3337GAT(1158)* ; 3386GAT(1186)
g1156 and 3336GAT(1169)* 3335GAT(1159)* ; 3383GAT(1187)
g1157 and 3334GAT(1171)* 3333GAT(1160)* ; 3380GAT(1188)
g1158 and 3332GAT(1172)* 3331GAT(1162)* ; 3377GAT(1189)
g1159 and 1044GAT(120)* 3344GAT(1163)* ; 3397GAT(1190)
g1160 and 3330GAT(1173)* 3329GAT(1164)* ; 3374GAT(1191)
g1161 and 996GAT(136)* 3341GAT(1156)* ; 3392GAT(1192)
g1162 and 3328GAT(1174)* 3327GAT(1166)* ; 3371GAT(1193)
g1163 and 3326GAT(1175)* 3325GAT(1168)* ; 3368GAT(1194)
g1164 and 3324GAT(1176)* 3323GAT(1170)* ; 3365GAT(1195)
g1165 and 3413GAT(1185)* 3260GAT(1109)* ; 3476GAT(1196)
g1166 and 3413GAT(1185)* 3362GAT(1149)* ; 3474GAT(1197)
g1167 and 3409GAT(1179)* 3408GAT(1178)* ; 3467GAT(1198)
g1168 and 3404GAT(1180)* 3353GAT(1153)* ; 3465GAT(1199)
g1169 and 3350GAT(1154)* 3404GAT(1180)* ; 3466GAT(1200)
g1170 and 3398GAT(1182)* 3401GAT(1181)* ; 3461GAT(1201)
g1171 and 3397GAT(1190)* 3396GAT(1183)* ; 3458GAT(1202)
g1172 and 3392GAT(1192)* 3239GAT(1116)* ; 3455GAT(1203)
g1173 and 3392GAT(1192)* 3341GAT(1156)* ; 3453GAT(1204)
g1174 and 1239GAT(55)* 3413GAT(1185)* ; 3475GAT(1205)
g1175 and 1191GAT(71)* 3410GAT(1177)* ; 3470GAT(1206)
g1176 and 996GAT(136)* 3392GAT(1192)* ; 3454GAT(1207)
g1177 and 948GAT(152)* 3389GAT(1184)* ; 3449GAT(1208)
g1178 and 900GAT(168)* 3386GAT(1186)* ; 3445GAT(1209)
g1179 and 852GAT(184)* 3383GAT(1187)* ; 3441GAT(1210)
g1180 and 804GAT(200)* 3380GAT(1188)* ; 3437GAT(1211)
g1181 and 756GAT(216)* 3377GAT(1189)* ; 3433GAT(1212)
g1182 and 708GAT(232)* 3374GAT(1191)* ; 3429GAT(1213)
g1183 and 660GAT(248)* 3371GAT(1193)* ; 3425GAT(1214)
g1184 and 612GAT(264)* 3368GAT(1194)* ; 3421GAT(1215)
g1185 and 564GAT(280)* 3365GAT(1195)* ; 3417GAT(1216)
g1186 and 3476GAT(1196)* 1287GAT(39)* ; 3548GAT(1217)
g1187 and 3475GAT(1205)* 3474GAT(1197)* ; 3545GAT(1218)
g1188 and 3470GAT(1206)* 3317GAT(1131)* ; 3542GAT(1219)
g1189 and 3470GAT(1206)* 3410GAT(1177)* ; 3540GAT(1220)
g1190 and 3466GAT(1200)* 3465GAT(1199)* ; 3533GAT(1221)
g1191 and 3461GAT(1201)* 3401GAT(1181)* ; 3531GAT(1222)
g1192 and 3398GAT(1182)* 3461GAT(1201)* ; 3532GAT(1223)
g1193 and 3455GAT(1203)* 3458GAT(1202)* ; 3527GAT(1224)
g1194 and 3454GAT(1207)* 3453GAT(1204)* ; 3524GAT(1225)
g1195 and 3449GAT(1208)* 3389GAT(1184)* ; 3519GAT(1226)
g1196 and 3445GAT(1209)* 3386GAT(1186)* ; 3514GAT(1227)
g1197 and 1191GAT(71)* 3470GAT(1206)* ; 3541GAT(1228)
g1198 and 3441GAT(1210)* 3383GAT(1187)* ; 3509GAT(1229)
g1199 and 1143GAT(87)* 3467GAT(1198)* ; 3536GAT(1230)
g1200 and 3437GAT(1211)* 3380GAT(1188)* ; 3504GAT(1231)
g1201 and 3433GAT(1212)* 3377GAT(1189)* ; 3499GAT(1232)
g1202 and 3429GAT(1213)* 3374GAT(1191)* ; 3494GAT(1233)
g1203 and 3449GAT(1208)* 3296GAT(1140)* ; 3521GAT(1234)
g1204 and 3425GAT(1214)* 3371GAT(1193)* ; 3489GAT(1235)
g1205 and 948GAT(152)* 3449GAT(1208)* ; 3520GAT(1236)
g1206 and 3445GAT(1209)* 3292GAT(1141)* ; 3516GAT(1237)
g1207 and 3421GAT(1215)* 3368GAT(1194)* ; 3484GAT(1238)
g1208 and 900GAT(168)* 3445GAT(1209)* ; 3515GAT(1239)
g1209 and 3441GAT(1210)* 3288GAT(1142)* ; 3511GAT(1240)
g1210 and 3417GAT(1216)* 3365GAT(1195)* ; 3479GAT(1241)
g1211 and 852GAT(184)* 3441GAT(1210)* ; 3510GAT(1242)
g1212 and 3437GAT(1211)* 3284GAT(1143)* ; 3506GAT(1243)
g1213 and 804GAT(200)* 3437GAT(1211)* ; 3505GAT(1244)
g1214 and 3433GAT(1212)* 3280GAT(1144)* ; 3501GAT(1245)
g1215 and 756GAT(216)* 3433GAT(1212)* ; 3500GAT(1246)
g1216 and 3429GAT(1213)* 3276GAT(1145)* ; 3496GAT(1247)
g1217 and 708GAT(232)* 3429GAT(1213)* ; 3495GAT(1248)
g1218 and 3425GAT(1214)* 3272GAT(1146)* ; 3491GAT(1249)
g1219 and 660GAT(248)* 3425GAT(1214)* ; 3490GAT(1250)
g1220 and 3421GAT(1215)* 3268GAT(1147)* ; 3486GAT(1251)
g1221 and 612GAT(264)* 3421GAT(1215)* ; 3485GAT(1252)
g1222 and 3417GAT(1216)* 3264GAT(1148)* ; 3481GAT(1253)
g1223 and 564GAT(280)* 3417GAT(1216)* ; 3480GAT(1254)
g1224 and 3548GAT(1217)* 1287GAT(39)* ; 3602GAT(1255)
g1225 and 3476GAT(1196)* 3548GAT(1217)* ; 3603GAT(1256)
g1226 and 3542GAT(1219)* 3545GAT(1218)* ; 3598GAT(1257)
g1227 and 3541GAT(1228)* 3540GAT(1220)* ; 3595GAT(1258)
g1228 and 3536GAT(1230)* 3356GAT(1152)* ; 3592GAT(1259)
g1229 and 3536GAT(1230)* 3467GAT(1198)* ; 3590GAT(1260)
g1230 and 3532GAT(1223)* 3531GAT(1222)* ; 3583GAT(1261)
g1231 and 3527GAT(1224)* 3458GAT(1202)* ; 3581GAT(1262)
g1232 and 3455GAT(1203)* 3527GAT(1224)* ; 3582GAT(1263)
g1233 and 3521GAT(1234)* 3524GAT(1225)* ; 3577GAT(1264)
g1234 and 3520GAT(1236)* 3519GAT(1226)* ; 3574GAT(1265)
g1235 and 3515GAT(1239)* 3514GAT(1227)* ; 3571GAT(1266)
g1236 and 3510GAT(1242)* 3509GAT(1229)* ; 3568GAT(1267)
g1237 and 1143GAT(87)* 3536GAT(1230)* ; 3591GAT(1268)
g1238 and 3505GAT(1244)* 3504GAT(1231)* ; 3565GAT(1269)
g1239 and 1095GAT(103)* 3533GAT(1221)* ; 3586GAT(1270)
g1240 and 3500GAT(1246)* 3499GAT(1232)* ; 3562GAT(1271)
g1241 and 3495GAT(1248)* 3494GAT(1233)* ; 3559GAT(1272)
g1242 and 3490GAT(1250)* 3489GAT(1235)* ; 3556GAT(1273)
g1243 and 3485GAT(1252)* 3484GAT(1238)* ; 3553GAT(1274)
g1244 and 3480GAT(1254)* 3479GAT(1241)* ; 3552GAT(1275)
g1245 and 3603GAT(1256)* 3602GAT(1255)* ; 3659GAT(1276)
g1246 and 3598GAT(1257)* 3545GAT(1218)* ; 3657GAT(1277)
g1247 and 3542GAT(1219)* 3598GAT(1257)* ; 3658GAT(1278)
g1248 and 3592GAT(1259)* 3595GAT(1258)* ; 3653GAT(1279)
g1249 and 3591GAT(1268)* 3590GAT(1260)* ; 3650GAT(1280)
g1250 and 3586GAT(1270)* 3404GAT(1180)* ; 3647GAT(1281)
g1251 and 3586GAT(1270)* 3533GAT(1221)* ; 3645GAT(1282)
g1252 and 3582GAT(1263)* 3581GAT(1262)* ; 3638GAT(1283)
g1253 and 3577GAT(1264)* 3524GAT(1225)* ; 3636GAT(1284)
g1254 and 1095GAT(103)* 3586GAT(1270)* ; 3646GAT(1285)
g1255 and 1047GAT(119)* 3583GAT(1261)* ; 3641GAT(1286)
g1256 and 3521GAT(1234)* 3577GAT(1264)* ; 3637GAT(1287)
g1257 and 3516GAT(1237)* 3574GAT(1265)* ; 3632GAT(1288)
g1258 and 3511GAT(1240)* 3571GAT(1266)* ; 3628GAT(1289)
g1259 and 3506GAT(1243)* 3568GAT(1267)* ; 3624GAT(1290)
g1260 and 3501GAT(1245)* 3565GAT(1269)* ; 3620GAT(1291)
g1261 and 3496GAT(1247)* 3562GAT(1271)* ; 3616GAT(1292)
g1262 and 3491GAT(1249)* 3559GAT(1272)* ; 3612GAT(1293)
g1263 and 3486GAT(1251)* 3556GAT(1273)* ; 3608GAT(1294)
g1264 and 3481GAT(1253)* 3553GAT(1274)* ; 3604GAT(1295)
g1265 and 3658GAT(1278)* 3657GAT(1277)* ; 3699GAT(1296)
g1266 and 3653GAT(1279)* 3595GAT(1258)* ; 3697GAT(1297)
g1267 and 3592GAT(1259)* 3653GAT(1279)* ; 3698GAT(1298)
g1268 and 3647GAT(1281)* 3650GAT(1280)* ; 3693GAT(1299)
g1269 and 3646GAT(1285)* 3645GAT(1282)* ; 3690GAT(1300)
g1270 and 3641GAT(1286)* 3461GAT(1201)* ; 3687GAT(1301)
g1271 and 3641GAT(1286)* 3583GAT(1261)* ; 3685GAT(1302)
g1272 and 3637GAT(1287)* 3636GAT(1284)* ; 3678GAT(1303)
g1273 and 3632GAT(1288)* 3574GAT(1265)* ; 3676GAT(1304)
g1274 and 1242GAT(54)* 3659GAT(1276)* ; 3702GAT(1305)
g1275 and 3628GAT(1289)* 3571GAT(1266)* ; 3674GAT(1306)
g1276 and 3624GAT(1290)* 3568GAT(1267)* ; 3672GAT(1307)
g1277 and 3620GAT(1291)* 3565GAT(1269)* ; 3670GAT(1308)
g1278 and 3616GAT(1292)* 3562GAT(1271)* ; 3668GAT(1309)
g1279 and 1047GAT(119)* 3641GAT(1286)* ; 3686GAT(1310)
g1280 and 3612GAT(1293)* 3559GAT(1272)* ; 3666GAT(1311)
g1281 and 999GAT(135)* 3638GAT(1283)* ; 3681GAT(1312)
g1282 and 3608GAT(1294)* 3556GAT(1273)* ; 3664GAT(1313)
g1283 and 3516GAT(1237)* 3632GAT(1288)* ; 3677GAT(1314)
g1284 and 3604GAT(1295)* 3553GAT(1274)* ; 3662GAT(1315)
g1285 and 3511GAT(1240)* 3628GAT(1289)* ; 3675GAT(1316)
g1286 and 3506GAT(1243)* 3624GAT(1290)* ; 3673GAT(1317)
g1287 and 3501GAT(1245)* 3620GAT(1291)* ; 3671GAT(1318)
g1288 and 3496GAT(1247)* 3616GAT(1292)* ; 3669GAT(1319)
g1289 and 3491GAT(1249)* 3612GAT(1293)* ; 3667GAT(1320)
g1290 and 3486GAT(1251)* 3608GAT(1294)* ; 3665GAT(1321)
g1291 and 3481GAT(1253)* 3604GAT(1295)* ; 3663GAT(1322)
g1292 and 3702GAT(1305)* 3548GAT(1217)* ; 3757GAT(1323)
g1293 and 3702GAT(1305)* 3659GAT(1276)* ; 3755GAT(1324)
g1294 and 3698GAT(1298)* 3697GAT(1297)* ; 3748GAT(1325)
g1295 and 3693GAT(1299)* 3650GAT(1280)* ; 3746GAT(1326)
g1296 and 3647GAT(1281)* 3693GAT(1299)* ; 3747GAT(1327)
g1297 and 3687GAT(1301)* 3690GAT(1300)* ; 3742GAT(1328)
g1298 and 3686GAT(1310)* 3685GAT(1302)* ; 3739GAT(1329)
g1299 and 3681GAT(1312)* 3527GAT(1224)* ; 3736GAT(1330)
g1300 and 3681GAT(1312)* 3638GAT(1283)* ; 3734GAT(1331)
g1301 and 3677GAT(1314)* 3676GAT(1304)* ; 3727GAT(1332)
g1302 and 1242GAT(54)* 3702GAT(1305)* ; 3756GAT(1333)
g1303 and 3675GAT(1316)* 3674GAT(1306)* ; 3724GAT(1334)
g1304 and 1194GAT(70)* 3699GAT(1296)* ; 3751GAT(1335)
g1305 and 3673GAT(1317)* 3672GAT(1307)* ; 3721GAT(1336)
g1306 and 3671GAT(1318)* 3670GAT(1308)* ; 3718GAT(1337)
g1307 and 3669GAT(1319)* 3668GAT(1309)* ; 3715GAT(1338)
g1308 and 3667GAT(1320)* 3666GAT(1311)* ; 3712GAT(1339)
g1309 and 999GAT(135)* 3681GAT(1312)* ; 3735GAT(1340)
g1310 and 3665GAT(1321)* 3664GAT(1313)* ; 3709GAT(1341)
g1311 and 951GAT(151)* 3678GAT(1303)* ; 3730GAT(1342)
g1312 and 3663GAT(1322)* 3662GAT(1315)* ; 3706GAT(1343)
g1313 and 3757GAT(1323)* 1290GAT(38)* ; 3821GAT(1344)
g1314 and 3756GAT(1333)* 3755GAT(1324)* ; 3818GAT(1345)
g1315 and 3751GAT(1335)* 3598GAT(1257)* ; 3815GAT(1346)
g1316 and 3751GAT(1335)* 3699GAT(1296)* ; 3813GAT(1347)
g1317 and 3747GAT(1327)* 3746GAT(1326)* ; 3806GAT(1348)
g1318 and 3742GAT(1328)* 3690GAT(1300)* ; 3804GAT(1349)
g1319 and 3687GAT(1301)* 3742GAT(1328)* ; 3805GAT(1350)
g1320 and 3736GAT(1330)* 3739GAT(1329)* ; 3800GAT(1351)
g1321 and 3735GAT(1340)* 3734GAT(1331)* ; 3797GAT(1352)
g1322 and 3730GAT(1342)* 3577GAT(1264)* ; 3794GAT(1353)
g1323 and 3730GAT(1342)* 3678GAT(1303)* ; 3792GAT(1354)
g1324 and 1194GAT(70)* 3751GAT(1335)* ; 3814GAT(1355)
g1325 and 1146GAT(86)* 3748GAT(1325)* ; 3809GAT(1356)
g1326 and 951GAT(151)* 3730GAT(1342)* ; 3793GAT(1357)
g1327 and 903GAT(167)* 3727GAT(1332)* ; 3788GAT(1358)
g1328 and 855GAT(183)* 3724GAT(1334)* ; 3784GAT(1359)
g1329 and 807GAT(199)* 3721GAT(1336)* ; 3780GAT(1360)
g1330 and 759GAT(215)* 3718GAT(1337)* ; 3776GAT(1361)
g1331 and 711GAT(231)* 3715GAT(1338)* ; 3772GAT(1362)
g1332 and 663GAT(247)* 3712GAT(1339)* ; 3768GAT(1363)
g1333 and 615GAT(263)* 3709GAT(1341)* ; 3764GAT(1364)
g1334 and 567GAT(279)* 3706GAT(1343)* ; 3760GAT(1365)
g1335 and 3821GAT(1344)* 1290GAT(38)* ; 3893GAT(1366)
g1336 and 3757GAT(1323)* 3821GAT(1344)* ; 3894GAT(1367)
g1337 and 3815GAT(1346)* 3818GAT(1345)* ; 3889GAT(1368)
g1338 and 3814GAT(1355)* 3813GAT(1347)* ; 3886GAT(1369)
g1339 and 3809GAT(1356)* 3653GAT(1279)* ; 3883GAT(1370)
g1340 and 3809GAT(1356)* 3748GAT(1325)* ; 3881GAT(1371)
g1341 and 3805GAT(1350)* 3804GAT(1349)* ; 3874GAT(1372)
g1342 and 3800GAT(1351)* 3739GAT(1329)* ; 3872GAT(1373)
g1343 and 3736GAT(1330)* 3800GAT(1351)* ; 3873GAT(1374)
g1344 and 3794GAT(1353)* 3797GAT(1352)* ; 3868GAT(1375)
g1345 and 3793GAT(1357)* 3792GAT(1354)* ; 3865GAT(1376)
g1346 and 3788GAT(1358)* 3727GAT(1332)* ; 3860GAT(1377)
g1347 and 3784GAT(1359)* 3724GAT(1334)* ; 3855GAT(1378)
g1348 and 3780GAT(1360)* 3721GAT(1336)* ; 3850GAT(1379)
g1349 and 1146GAT(86)* 3809GAT(1356)* ; 3882GAT(1380)
g1350 and 3776GAT(1361)* 3718GAT(1337)* ; 3845GAT(1381)
g1351 and 1098GAT(102)* 3806GAT(1348)* ; 3877GAT(1382)
g1352 and 3772GAT(1362)* 3715GAT(1338)* ; 3840GAT(1383)
g1353 and 3768GAT(1363)* 3712GAT(1339)* ; 3835GAT(1384)
g1354 and 3764GAT(1364)* 3709GAT(1341)* ; 3830GAT(1385)
g1355 and 3788GAT(1358)* 3632GAT(1288)* ; 3862GAT(1386)
g1356 and 3760GAT(1365)* 3706GAT(1343)* ; 3825GAT(1387)
g1357 and 903GAT(167)* 3788GAT(1358)* ; 3861GAT(1388)
g1358 and 3784GAT(1359)* 3628GAT(1289)* ; 3857GAT(1389)
g1359 and 855GAT(183)* 3784GAT(1359)* ; 3856GAT(1390)
g1360 and 3780GAT(1360)* 3624GAT(1290)* ; 3852GAT(1391)
g1361 and 807GAT(199)* 3780GAT(1360)* ; 3851GAT(1392)
g1362 and 3776GAT(1361)* 3620GAT(1291)* ; 3847GAT(1393)
g1363 and 759GAT(215)* 3776GAT(1361)* ; 3846GAT(1394)
g1364 and 3772GAT(1362)* 3616GAT(1292)* ; 3842GAT(1395)
g1365 and 711GAT(231)* 3772GAT(1362)* ; 3841GAT(1396)
g1366 and 3768GAT(1363)* 3612GAT(1293)* ; 3837GAT(1397)
g1367 and 663GAT(247)* 3768GAT(1363)* ; 3836GAT(1398)
g1368 and 3764GAT(1364)* 3608GAT(1294)* ; 3832GAT(1399)
g1369 and 615GAT(263)* 3764GAT(1364)* ; 3831GAT(1400)
g1370 and 3760GAT(1365)* 3604GAT(1295)* ; 3827GAT(1401)
g1371 and 567GAT(279)* 3760GAT(1365)* ; 3826GAT(1402)
g1372 and 3894GAT(1367)* 3893GAT(1366)* ; 3944GAT(1403)
g1373 and 3889GAT(1368)* 3818GAT(1345)* ; 3942GAT(1404)
g1374 and 3815GAT(1346)* 3889GAT(1368)* ; 3943GAT(1405)
g1375 and 3883GAT(1370)* 3886GAT(1369)* ; 3938GAT(1406)
g1376 and 3882GAT(1380)* 3881GAT(1371)* ; 3935GAT(1407)
g1377 and 3877GAT(1382)* 3693GAT(1299)* ; 3932GAT(1408)
g1378 and 3877GAT(1382)* 3806GAT(1348)* ; 3930GAT(1409)
g1379 and 3873GAT(1374)* 3872GAT(1373)* ; 3923GAT(1410)
g1380 and 3868GAT(1375)* 3797GAT(1352)* ; 3921GAT(1411)
g1381 and 3794GAT(1353)* 3868GAT(1375)* ; 3922GAT(1412)
g1382 and 3862GAT(1386)* 3865GAT(1376)* ; 3917GAT(1413)
g1383 and 3861GAT(1388)* 3860GAT(1377)* ; 3914GAT(1414)
g1384 and 3856GAT(1390)* 3855GAT(1378)* ; 3911GAT(1415)
g1385 and 3851GAT(1392)* 3850GAT(1379)* ; 3908GAT(1416)
g1386 and 3846GAT(1394)* 3845GAT(1381)* ; 3905GAT(1417)
g1387 and 1098GAT(102)* 3877GAT(1382)* ; 3931GAT(1418)
g1388 and 3841GAT(1396)* 3840GAT(1383)* ; 3902GAT(1419)
g1389 and 1050GAT(118)* 3874GAT(1372)* ; 3926GAT(1420)
g1390 and 3836GAT(1398)* 3835GAT(1384)* ; 3899GAT(1421)
g1391 and 3831GAT(1400)* 3830GAT(1385)* ; 3896GAT(1422)
g1392 and 3826GAT(1402)* 3825GAT(1387)* ; 3895GAT(1423)
g1393 and 3943GAT(1405)* 3942GAT(1404)* ; 3998GAT(1424)
g1394 and 3938GAT(1406)* 3886GAT(1369)* ; 3996GAT(1425)
g1395 and 3883GAT(1370)* 3938GAT(1406)* ; 3997GAT(1426)
g1396 and 3932GAT(1408)* 3935GAT(1407)* ; 3992GAT(1427)
g1397 and 3931GAT(1418)* 3930GAT(1409)* ; 3989GAT(1428)
g1398 and 3926GAT(1420)* 3742GAT(1328)* ; 3986GAT(1429)
g1399 and 3926GAT(1420)* 3874GAT(1372)* ; 3984GAT(1430)
g1400 and 3922GAT(1412)* 3921GAT(1411)* ; 3977GAT(1431)
g1401 and 3917GAT(1413)* 3865GAT(1376)* ; 3975GAT(1432)
g1402 and 1245GAT(53)* 3944GAT(1403)* ; 4001GAT(1433)
g1403 and 1050GAT(118)* 3926GAT(1420)* ; 3985GAT(1434)
g1404 and 1002GAT(134)* 3923GAT(1410)* ; 3980GAT(1435)
g1405 and 3862GAT(1386)* 3917GAT(1413)* ; 3976GAT(1436)
g1406 and 3857GAT(1389)* 3914GAT(1414)* ; 3971GAT(1437)
g1407 and 3852GAT(1391)* 3911GAT(1415)* ; 3967GAT(1438)
g1408 and 3847GAT(1393)* 3908GAT(1416)* ; 3963GAT(1439)
g1409 and 3842GAT(1395)* 3905GAT(1417)* ; 3959GAT(1440)
g1410 and 3837GAT(1397)* 3902GAT(1419)* ; 3955GAT(1441)
g1411 and 3832GAT(1399)* 3899GAT(1421)* ; 3951GAT(1442)
g1412 and 3827GAT(1401)* 3896GAT(1422)* ; 3947GAT(1443)
g1413 and 4001GAT(1433)* 3821GAT(1344)* ; 4049GAT(1444)
g1414 and 4001GAT(1433)* 3944GAT(1403)* ; 4047GAT(1445)
g1415 and 3997GAT(1426)* 3996GAT(1425)* ; 4040GAT(1446)
g1416 and 3992GAT(1427)* 3935GAT(1407)* ; 4038GAT(1447)
g1417 and 3932GAT(1408)* 3992GAT(1427)* ; 4039GAT(1448)
g1418 and 3986GAT(1429)* 3989GAT(1428)* ; 4034GAT(1449)
g1419 and 3985GAT(1434)* 3984GAT(1430)* ; 4031GAT(1450)
g1420 and 3980GAT(1435)* 3800GAT(1351)* ; 4028GAT(1451)
g1421 and 3980GAT(1435)* 3923GAT(1410)* ; 4026GAT(1452)
g1422 and 3976GAT(1436)* 3975GAT(1432)* ; 4019GAT(1453)
g1423 and 3971GAT(1437)* 3914GAT(1414)* ; 4017GAT(1454)
g1424 and 1245GAT(53)* 4001GAT(1433)* ; 4048GAT(1455)
g1425 and 3967GAT(1438)* 3911GAT(1415)* ; 4015GAT(1456)
g1426 and 1197GAT(69)* 3998GAT(1424)* ; 4043GAT(1457)
g1427 and 3963GAT(1439)* 3908GAT(1416)* ; 4013GAT(1458)
g1428 and 3959GAT(1440)* 3905GAT(1417)* ; 4011GAT(1459)
g1429 and 3955GAT(1441)* 3902GAT(1419)* ; 4009GAT(1460)
g1430 and 3951GAT(1442)* 3899GAT(1421)* ; 4007GAT(1461)
g1431 and 1002GAT(134)* 3980GAT(1435)* ; 4027GAT(1462)
g1432 and 3947GAT(1443)* 3896GAT(1422)* ; 4005GAT(1463)
g1433 and 954GAT(150)* 3977GAT(1431)* ; 4022GAT(1464)
g1434 and 3857GAT(1389)* 3971GAT(1437)* ; 4018GAT(1465)
g1435 and 3852GAT(1391)* 3967GAT(1438)* ; 4016GAT(1466)
g1436 and 3847GAT(1393)* 3963GAT(1439)* ; 4014GAT(1467)
g1437 and 3842GAT(1395)* 3959GAT(1440)* ; 4012GAT(1468)
g1438 and 3837GAT(1397)* 3955GAT(1441)* ; 4010GAT(1469)
g1439 and 3832GAT(1399)* 3951GAT(1442)* ; 4008GAT(1470)
g1440 and 3827GAT(1401)* 3947GAT(1443)* ; 4006GAT(1471)
g1441 and 4049GAT(1444)* 1293GAT(37)* ; 4106GAT(1472)
g1442 and 4048GAT(1455)* 4047GAT(1445)* ; 4103GAT(1473)
g1443 and 4043GAT(1457)* 3889GAT(1368)* ; 4100GAT(1474)
g1444 and 4043GAT(1457)* 3998GAT(1424)* ; 4098GAT(1475)
g1445 and 4039GAT(1448)* 4038GAT(1447)* ; 4091GAT(1476)
g1446 and 4034GAT(1449)* 3989GAT(1428)* ; 4089GAT(1477)
g1447 and 3986GAT(1429)* 4034GAT(1449)* ; 4090GAT(1478)
g1448 and 4028GAT(1451)* 4031GAT(1450)* ; 4085GAT(1479)
g1449 and 4027GAT(1462)* 4026GAT(1452)* ; 4082GAT(1480)
g1450 and 4022GAT(1464)* 3868GAT(1375)* ; 4079GAT(1481)
g1451 and 4022GAT(1464)* 3977GAT(1431)* ; 4077GAT(1482)
g1452 and 4018GAT(1465)* 4017GAT(1454)* ; 4070GAT(1483)
g1453 and 4016GAT(1466)* 4015GAT(1456)* ; 4067GAT(1484)
g1454 and 1197GAT(69)* 4043GAT(1457)* ; 4099GAT(1485)
g1455 and 4014GAT(1467)* 4013GAT(1458)* ; 4064GAT(1486)
g1456 and 1149GAT(85)* 4040GAT(1446)* ; 4094GAT(1487)
g1457 and 4012GAT(1468)* 4011GAT(1459)* ; 4061GAT(1488)
g1458 and 4010GAT(1469)* 4009GAT(1460)* ; 4058GAT(1489)
g1459 and 4008GAT(1470)* 4007GAT(1461)* ; 4055GAT(1490)
g1460 and 4006GAT(1471)* 4005GAT(1463)* ; 4052GAT(1491)
g1461 and 954GAT(150)* 4022GAT(1464)* ; 4078GAT(1492)
g1462 and 906GAT(166)* 4019GAT(1453)* ; 4073GAT(1493)
g1463 and 4106GAT(1472)* 1293GAT(37)* ; 4171GAT(1494)
g1464 and 4049GAT(1444)* 4106GAT(1472)* ; 4172GAT(1495)
g1465 and 4100GAT(1474)* 4103GAT(1473)* ; 4167GAT(1496)
g1466 and 4099GAT(1485)* 4098GAT(1475)* ; 4164GAT(1497)
g1467 and 4094GAT(1487)* 3938GAT(1406)* ; 4161GAT(1498)
g1468 and 4094GAT(1487)* 4040GAT(1446)* ; 4159GAT(1499)
g1469 and 4090GAT(1478)* 4089GAT(1477)* ; 4152GAT(1500)
g1470 and 4085GAT(1479)* 4031GAT(1450)* ; 4150GAT(1501)
g1471 and 4028GAT(1451)* 4085GAT(1479)* ; 4151GAT(1502)
g1472 and 4079GAT(1481)* 4082GAT(1480)* ; 4146GAT(1503)
g1473 and 4078GAT(1492)* 4077GAT(1482)* ; 4143GAT(1504)
g1474 and 4073GAT(1493)* 3917GAT(1413)* ; 4140GAT(1505)
g1475 and 4073GAT(1493)* 4019GAT(1453)* ; 4138GAT(1506)
g1476 and 1149GAT(85)* 4094GAT(1487)* ; 4160GAT(1507)
g1477 and 1101GAT(101)* 4091GAT(1476)* ; 4155GAT(1508)
g1478 and 906GAT(166)* 4073GAT(1493)* ; 4139GAT(1509)
g1479 and 858GAT(182)* 4070GAT(1483)* ; 4134GAT(1510)
g1480 and 810GAT(198)* 4067GAT(1484)* ; 4130GAT(1511)
g1481 and 762GAT(214)* 4064GAT(1486)* ; 4126GAT(1512)
g1482 and 714GAT(230)* 4061GAT(1488)* ; 4122GAT(1513)
g1483 and 666GAT(246)* 4058GAT(1489)* ; 4118GAT(1514)
g1484 and 618GAT(262)* 4055GAT(1490)* ; 4114GAT(1515)
g1485 and 570GAT(278)* 4052GAT(1491)* ; 4110GAT(1516)
g1486 and 4172GAT(1495)* 4171GAT(1494)* ; 4238GAT(1517)
g1487 and 4167GAT(1496)* 4103GAT(1473)* ; 4236GAT(1518)
g1488 and 4100GAT(1474)* 4167GAT(1496)* ; 4237GAT(1519)
g1489 and 4161GAT(1498)* 4164GAT(1497)* ; 4232GAT(1520)
g1490 and 4160GAT(1507)* 4159GAT(1499)* ; 4229GAT(1521)
g1491 and 4155GAT(1508)* 3992GAT(1427)* ; 4226GAT(1522)
g1492 and 4155GAT(1508)* 4091GAT(1476)* ; 4224GAT(1523)
g1493 and 4151GAT(1502)* 4150GAT(1501)* ; 4217GAT(1524)
g1494 and 4146GAT(1503)* 4082GAT(1480)* ; 4215GAT(1525)
g1495 and 4079GAT(1481)* 4146GAT(1503)* ; 4216GAT(1526)
g1496 and 4140GAT(1505)* 4143GAT(1504)* ; 4211GAT(1527)
g1497 and 4139GAT(1509)* 4138GAT(1506)* ; 4208GAT(1528)
g1498 and 4134GAT(1510)* 4070GAT(1483)* ; 4203GAT(1529)
g1499 and 4130GAT(1511)* 4067GAT(1484)* ; 4198GAT(1530)
g1500 and 4126GAT(1512)* 4064GAT(1486)* ; 4193GAT(1531)
g1501 and 4122GAT(1513)* 4061GAT(1488)* ; 4188GAT(1532)
g1502 and 1101GAT(101)* 4155GAT(1508)* ; 4225GAT(1533)
g1503 and 4118GAT(1514)* 4058GAT(1489)* ; 4183GAT(1534)
g1504 and 1053GAT(117)* 4152GAT(1500)* ; 4220GAT(1535)
g1505 and 4114GAT(1515)* 4055GAT(1490)* ; 4178GAT(1536)
g1506 and 4110GAT(1516)* 4052GAT(1491)* ; 4173GAT(1537)
g1507 and 4134GAT(1510)* 3971GAT(1437)* ; 4205GAT(1538)
g1508 and 858GAT(182)* 4134GAT(1510)* ; 4204GAT(1539)
g1509 and 4130GAT(1511)* 3967GAT(1438)* ; 4200GAT(1540)
g1510 and 810GAT(198)* 4130GAT(1511)* ; 4199GAT(1541)
g1511 and 4126GAT(1512)* 3963GAT(1439)* ; 4195GAT(1542)
g1512 and 762GAT(214)* 4126GAT(1512)* ; 4194GAT(1543)
g1513 and 4122GAT(1513)* 3959GAT(1440)* ; 4190GAT(1544)
g1514 and 714GAT(230)* 4122GAT(1513)* ; 4189GAT(1545)
g1515 and 4118GAT(1514)* 3955GAT(1441)* ; 4185GAT(1546)
g1516 and 666GAT(246)* 4118GAT(1514)* ; 4184GAT(1547)
g1517 and 4114GAT(1515)* 3951GAT(1442)* ; 4180GAT(1548)
g1518 and 618GAT(262)* 4114GAT(1515)* ; 4179GAT(1549)
g1519 and 4110GAT(1516)* 3947GAT(1443)* ; 4175GAT(1550)
g1520 and 570GAT(278)* 4110GAT(1516)* ; 4174GAT(1551)
g1521 and 4237GAT(1519)* 4236GAT(1518)* ; 4287GAT(1552)
g1522 and 4232GAT(1520)* 4164GAT(1497)* ; 4285GAT(1553)
g1523 and 4161GAT(1498)* 4232GAT(1520)* ; 4286GAT(1554)
g1524 and 4226GAT(1522)* 4229GAT(1521)* ; 4281GAT(1555)
g1525 and 4225GAT(1533)* 4224GAT(1523)* ; 4278GAT(1556)
g1526 and 4220GAT(1535)* 4034GAT(1449)* ; 4275GAT(1557)
g1527 and 4220GAT(1535)* 4152GAT(1500)* ; 4273GAT(1558)
g1528 and 4216GAT(1526)* 4215GAT(1525)* ; 4266GAT(1559)
g1529 and 4211GAT(1527)* 4143GAT(1504)* ; 4264GAT(1560)
g1530 and 4140GAT(1505)* 4211GAT(1527)* ; 4265GAT(1561)
g1531 and 4205GAT(1538)* 4208GAT(1528)* ; 4260GAT(1562)
g1532 and 4204GAT(1539)* 4203GAT(1529)* ; 4257GAT(1563)
g1533 and 1248GAT(52)* 4238GAT(1517)* ; 4290GAT(1564)
g1534 and 4199GAT(1541)* 4198GAT(1530)* ; 4254GAT(1565)
g1535 and 4194GAT(1543)* 4193GAT(1531)* ; 4251GAT(1566)
g1536 and 4189GAT(1545)* 4188GAT(1532)* ; 4248GAT(1567)
g1537 and 4184GAT(1547)* 4183GAT(1534)* ; 4245GAT(1568)
g1538 and 1053GAT(117)* 4220GAT(1535)* ; 4274GAT(1569)
g1539 and 4179GAT(1549)* 4178GAT(1536)* ; 4242GAT(1570)
g1540 and 1005GAT(133)* 4217GAT(1524)* ; 4269GAT(1571)
g1541 and 4174GAT(1551)* 4173GAT(1537)* ; 4241GAT(1572)
g1542 and 4290GAT(1564)* 4106GAT(1472)* ; 4350GAT(1573)
g1543 and 4290GAT(1564)* 4238GAT(1517)* ; 4348GAT(1574)
g1544 and 4286GAT(1554)* 4285GAT(1553)* ; 4341GAT(1575)
g1545 and 4281GAT(1555)* 4229GAT(1521)* ; 4339GAT(1576)
g1546 and 4226GAT(1522)* 4281GAT(1555)* ; 4340GAT(1577)
g1547 and 4275GAT(1557)* 4278GAT(1556)* ; 4335GAT(1578)
g1548 and 4274GAT(1569)* 4273GAT(1558)* ; 4332GAT(1579)
g1549 and 4269GAT(1571)* 4085GAT(1479)* ; 4329GAT(1580)
g1550 and 4269GAT(1571)* 4217GAT(1524)* ; 4327GAT(1581)
g1551 and 4265GAT(1561)* 4264GAT(1560)* ; 4320GAT(1582)
g1552 and 4260GAT(1562)* 4208GAT(1528)* ; 4318GAT(1583)
g1553 and 1248GAT(52)* 4290GAT(1564)* ; 4349GAT(1584)
g1554 and 1200GAT(68)* 4287GAT(1552)* ; 4344GAT(1585)
g1555 and 1005GAT(133)* 4269GAT(1571)* ; 4328GAT(1586)
g1556 and 957GAT(149)* 4266GAT(1559)* ; 4323GAT(1587)
g1557 and 4205GAT(1538)* 4260GAT(1562)* ; 4319GAT(1588)
g1558 and 4200GAT(1540)* 4257GAT(1563)* ; 4314GAT(1589)
g1559 and 4195GAT(1542)* 4254GAT(1565)* ; 4310GAT(1590)
g1560 and 4190GAT(1544)* 4251GAT(1566)* ; 4306GAT(1591)
g1561 and 4185GAT(1546)* 4248GAT(1567)* ; 4302GAT(1592)
g1562 and 4180GAT(1548)* 4245GAT(1568)* ; 4298GAT(1593)
g1563 and 4175GAT(1550)* 4242GAT(1570)* ; 4294GAT(1594)
g1564 and 4350GAT(1573)* 1296GAT(36)* ; 4401GAT(1595)
g1565 and 4349GAT(1584)* 4348GAT(1574)* ; 4398GAT(1596)
g1566 and 4344GAT(1585)* 4167GAT(1496)* ; 4395GAT(1597)
g1567 and 4344GAT(1585)* 4287GAT(1552)* ; 4393GAT(1598)
g1568 and 4340GAT(1577)* 4339GAT(1576)* ; 4386GAT(1599)
g1569 and 4335GAT(1578)* 4278GAT(1556)* ; 4384GAT(1600)
g1570 and 4275GAT(1557)* 4335GAT(1578)* ; 4385GAT(1601)
g1571 and 4329GAT(1580)* 4332GAT(1579)* ; 4380GAT(1602)
g1572 and 4328GAT(1586)* 4327GAT(1581)* ; 4377GAT(1603)
g1573 and 4323GAT(1587)* 4146GAT(1503)* ; 4374GAT(1604)
g1574 and 4323GAT(1587)* 4266GAT(1559)* ; 4372GAT(1605)
g1575 and 4319GAT(1588)* 4318GAT(1583)* ; 4365GAT(1606)
g1576 and 4314GAT(1589)* 4257GAT(1563)* ; 4363GAT(1607)
g1577 and 4310GAT(1590)* 4254GAT(1565)* ; 4361GAT(1608)
g1578 and 1200GAT(68)* 4344GAT(1585)* ; 4394GAT(1609)
g1579 and 4306GAT(1591)* 4251GAT(1566)* ; 4359GAT(1610)
g1580 and 1152GAT(84)* 4341GAT(1575)* ; 4389GAT(1611)
g1581 and 4302GAT(1592)* 4248GAT(1567)* ; 4357GAT(1612)
g1582 and 4298GAT(1593)* 4245GAT(1568)* ; 4355GAT(1613)
g1583 and 4294GAT(1594)* 4242GAT(1570)* ; 4353GAT(1614)
g1584 and 957GAT(149)* 4323GAT(1587)* ; 4373GAT(1615)
g1585 and 909GAT(165)* 4320GAT(1582)* ; 4368GAT(1616)
g1586 and 4200GAT(1540)* 4314GAT(1589)* ; 4364GAT(1617)
g1587 and 4195GAT(1542)* 4310GAT(1590)* ; 4362GAT(1618)
g1588 and 4190GAT(1544)* 4306GAT(1591)* ; 4360GAT(1619)
g1589 and 4185GAT(1546)* 4302GAT(1592)* ; 4358GAT(1620)
g1590 and 4180GAT(1548)* 4298GAT(1593)* ; 4356GAT(1621)
g1591 and 4175GAT(1550)* 4294GAT(1594)* ; 4354GAT(1622)
g1592 and 4401GAT(1595)* 1296GAT(36)* ; 4460GAT(1623)
g1593 and 4350GAT(1573)* 4401GAT(1595)* ; 4461GAT(1624)
g1594 and 4395GAT(1597)* 4398GAT(1596)* ; 4456GAT(1625)
g1595 and 4394GAT(1609)* 4393GAT(1598)* ; 4453GAT(1626)
g1596 and 4389GAT(1611)* 4232GAT(1520)* ; 4450GAT(1627)
g1597 and 4389GAT(1611)* 4341GAT(1575)* ; 4448GAT(1628)
g1598 and 4385GAT(1601)* 4384GAT(1600)* ; 4441GAT(1629)
g1599 and 4380GAT(1602)* 4332GAT(1579)* ; 4439GAT(1630)
g1600 and 4329GAT(1580)* 4380GAT(1602)* ; 4440GAT(1631)
g1601 and 4374GAT(1604)* 4377GAT(1603)* ; 4435GAT(1632)
g1602 and 4373GAT(1615)* 4372GAT(1605)* ; 4432GAT(1633)
g1603 and 4368GAT(1616)* 4211GAT(1527)* ; 4429GAT(1634)
g1604 and 4368GAT(1616)* 4320GAT(1582)* ; 4427GAT(1635)
g1605 and 4364GAT(1617)* 4363GAT(1607)* ; 4420GAT(1636)
g1606 and 4362GAT(1618)* 4361GAT(1608)* ; 4417GAT(1637)
g1607 and 4360GAT(1619)* 4359GAT(1610)* ; 4414GAT(1638)
g1608 and 1152GAT(84)* 4389GAT(1611)* ; 4449GAT(1639)
g1609 and 4358GAT(1620)* 4357GAT(1612)* ; 4411GAT(1640)
g1610 and 1104GAT(100)* 4386GAT(1599)* ; 4444GAT(1641)
g1611 and 4356GAT(1621)* 4355GAT(1613)* ; 4408GAT(1642)
g1612 and 4354GAT(1622)* 4353GAT(1614)* ; 4405GAT(1643)
g1613 and 909GAT(165)* 4368GAT(1616)* ; 4428GAT(1644)
g1614 and 861GAT(181)* 4365GAT(1606)* ; 4423GAT(1645)
g1615 and 4461GAT(1624)* 4460GAT(1623)* ; 4521GAT(1646)
g1616 and 4456GAT(1625)* 4398GAT(1596)* ; 4519GAT(1647)
g1617 and 4395GAT(1597)* 4456GAT(1625)* ; 4520GAT(1648)
g1618 and 4450GAT(1627)* 4453GAT(1626)* ; 4515GAT(1649)
g1619 and 4449GAT(1639)* 4448GAT(1628)* ; 4512GAT(1650)
g1620 and 4444GAT(1641)* 4281GAT(1555)* ; 4509GAT(1651)
g1621 and 4444GAT(1641)* 4386GAT(1599)* ; 4507GAT(1652)
g1622 and 4440GAT(1631)* 4439GAT(1630)* ; 4500GAT(1653)
g1623 and 4435GAT(1632)* 4377GAT(1603)* ; 4498GAT(1654)
g1624 and 4374GAT(1604)* 4435GAT(1632)* ; 4499GAT(1655)
g1625 and 4429GAT(1634)* 4432GAT(1633)* ; 4494GAT(1656)
g1626 and 4428GAT(1644)* 4427GAT(1635)* ; 4491GAT(1657)
g1627 and 4423GAT(1645)* 4260GAT(1562)* ; 4488GAT(1658)
g1628 and 4423GAT(1645)* 4365GAT(1606)* ; 4486GAT(1659)
g1629 and 1104GAT(100)* 4444GAT(1641)* ; 4508GAT(1660)
g1630 and 1056GAT(116)* 4441GAT(1629)* ; 4503GAT(1661)
g1631 and 861GAT(181)* 4423GAT(1645)* ; 4487GAT(1662)
g1632 and 813GAT(197)* 4420GAT(1636)* ; 4482GAT(1663)
g1633 and 765GAT(213)* 4417GAT(1637)* ; 4478GAT(1664)
g1634 and 717GAT(229)* 4414GAT(1638)* ; 4474GAT(1665)
g1635 and 669GAT(245)* 4411GAT(1640)* ; 4470GAT(1666)
g1636 and 621GAT(261)* 4408GAT(1642)* ; 4466GAT(1667)
g1637 and 573GAT(277)* 4405GAT(1643)* ; 4462GAT(1668)
g1638 and 4520GAT(1648)* 4519GAT(1647)* ; 4584GAT(1669)
g1639 and 4515GAT(1649)* 4453GAT(1626)* ; 4582GAT(1670)
g1640 and 4450GAT(1627)* 4515GAT(1649)* ; 4583GAT(1671)
g1641 and 4509GAT(1651)* 4512GAT(1650)* ; 4578GAT(1672)
g1642 and 4508GAT(1660)* 4507GAT(1652)* ; 4575GAT(1673)
g1643 and 4503GAT(1661)* 4335GAT(1578)* ; 4572GAT(1674)
g1644 and 4503GAT(1661)* 4441GAT(1629)* ; 4570GAT(1675)
g1645 and 4499GAT(1655)* 4498GAT(1654)* ; 4563GAT(1676)
g1646 and 4494GAT(1656)* 4432GAT(1633)* ; 4561GAT(1677)
g1647 and 4429GAT(1634)* 4494GAT(1656)* ; 4562GAT(1678)
g1648 and 4488GAT(1658)* 4491GAT(1657)* ; 4557GAT(1679)
g1649 and 4487GAT(1662)* 4486GAT(1659)* ; 4554GAT(1680)
g1650 and 4482GAT(1663)* 4420GAT(1636)* ; 4549GAT(1681)
g1651 and 1251GAT(51)* 4521GAT(1646)* ; 4587GAT(1682)
g1652 and 4478GAT(1664)* 4417GAT(1637)* ; 4544GAT(1683)
g1653 and 4474GAT(1665)* 4414GAT(1638)* ; 4539GAT(1684)
g1654 and 4470GAT(1666)* 4411GAT(1640)* ; 4534GAT(1685)
g1655 and 4466GAT(1667)* 4408GAT(1642)* ; 4529GAT(1686)
g1656 and 1056GAT(116)* 4503GAT(1661)* ; 4571GAT(1687)
g1657 and 4462GAT(1668)* 4405GAT(1643)* ; 4524GAT(1688)
g1658 and 1008GAT(132)* 4500GAT(1653)* ; 4566GAT(1689)
g1659 and 4482GAT(1663)* 4314GAT(1589)* ; 4551GAT(1690)
g1660 and 813GAT(197)* 4482GAT(1663)* ; 4550GAT(1691)
g1661 and 4478GAT(1664)* 4310GAT(1590)* ; 4546GAT(1692)
g1662 and 765GAT(213)* 4478GAT(1664)* ; 4545GAT(1693)
g1663 and 4474GAT(1665)* 4306GAT(1591)* ; 4541GAT(1694)
g1664 and 717GAT(229)* 4474GAT(1665)* ; 4540GAT(1695)
g1665 and 4470GAT(1666)* 4302GAT(1592)* ; 4536GAT(1696)
g1666 and 669GAT(245)* 4470GAT(1666)* ; 4535GAT(1697)
g1667 and 4466GAT(1667)* 4298GAT(1593)* ; 4531GAT(1698)
g1668 and 621GAT(261)* 4466GAT(1667)* ; 4530GAT(1699)
g1669 and 4462GAT(1668)* 4294GAT(1594)* ; 4526GAT(1700)
g1670 and 573GAT(277)* 4462GAT(1668)* ; 4525GAT(1701)
g1671 and 4587GAT(1682)* 4401GAT(1595)* ; 4643GAT(1702)
g1672 and 4587GAT(1682)* 4521GAT(1646)* ; 4641GAT(1703)
g1673 and 4583GAT(1671)* 4582GAT(1670)* ; 4634GAT(1704)
g1674 and 4578GAT(1672)* 4512GAT(1650)* ; 4632GAT(1705)
g1675 and 4509GAT(1651)* 4578GAT(1672)* ; 4633GAT(1706)
g1676 and 4572GAT(1674)* 4575GAT(1673)* ; 4628GAT(1707)
g1677 and 4571GAT(1687)* 4570GAT(1675)* ; 4625GAT(1708)
g1678 and 4566GAT(1689)* 4380GAT(1602)* ; 4622GAT(1709)
g1679 and 4566GAT(1689)* 4500GAT(1653)* ; 4620GAT(1710)
g1680 and 4562GAT(1678)* 4561GAT(1677)* ; 4613GAT(1711)
g1681 and 4557GAT(1679)* 4491GAT(1657)* ; 4611GAT(1712)
g1682 and 4488GAT(1658)* 4557GAT(1679)* ; 4612GAT(1713)
g1683 and 4551GAT(1690)* 4554GAT(1680)* ; 4607GAT(1714)
g1684 and 4550GAT(1691)* 4549GAT(1681)* ; 4604GAT(1715)
g1685 and 1251GAT(51)* 4587GAT(1682)* ; 4642GAT(1716)
g1686 and 4545GAT(1693)* 4544GAT(1683)* ; 4601GAT(1717)
g1687 and 1203GAT(67)* 4584GAT(1669)* ; 4637GAT(1718)
g1688 and 4540GAT(1695)* 4539GAT(1684)* ; 4598GAT(1719)
g1689 and 4535GAT(1697)* 4534GAT(1685)* ; 4595GAT(1720)
g1690 and 4530GAT(1699)* 4529GAT(1686)* ; 4592GAT(1721)
g1691 and 4525GAT(1701)* 4524GAT(1688)* ; 4591GAT(1722)
g1692 and 1008GAT(132)* 4566GAT(1689)* ; 4621GAT(1723)
g1693 and 960GAT(148)* 4563GAT(1676)* ; 4616GAT(1724)
g1694 and 4643GAT(1702)* 1299GAT(35)* ; 4704GAT(1725)
g1695 and 4642GAT(1716)* 4641GAT(1703)* ; 4701GAT(1726)
g1696 and 4637GAT(1718)* 4456GAT(1625)* ; 4698GAT(1727)
g1697 and 4637GAT(1718)* 4584GAT(1669)* ; 4696GAT(1728)
g1698 and 4633GAT(1706)* 4632GAT(1705)* ; 4689GAT(1729)
g1699 and 4628GAT(1707)* 4575GAT(1673)* ; 4687GAT(1730)
g1700 and 4572GAT(1674)* 4628GAT(1707)* ; 4688GAT(1731)
g1701 and 4622GAT(1709)* 4625GAT(1708)* ; 4683GAT(1732)
g1702 and 4621GAT(1723)* 4620GAT(1710)* ; 4680GAT(1733)
g1703 and 4616GAT(1724)* 4435GAT(1632)* ; 4677GAT(1734)
g1704 and 4616GAT(1724)* 4563GAT(1676)* ; 4675GAT(1735)
g1705 and 4612GAT(1713)* 4611GAT(1712)* ; 4668GAT(1736)
g1706 and 4607GAT(1714)* 4554GAT(1680)* ; 4666GAT(1737)
g1707 and 1203GAT(67)* 4637GAT(1718)* ; 4697GAT(1738)
g1708 and 1155GAT(83)* 4634GAT(1704)* ; 4692GAT(1739)
g1709 and 960GAT(148)* 4616GAT(1724)* ; 4676GAT(1740)
g1710 and 912GAT(164)* 4613GAT(1711)* ; 4671GAT(1741)
g1711 and 4551GAT(1690)* 4607GAT(1714)* ; 4667GAT(1742)
g1712 and 4546GAT(1692)* 4604GAT(1715)* ; 4662GAT(1743)
g1713 and 4541GAT(1694)* 4601GAT(1717)* ; 4658GAT(1744)
g1714 and 4536GAT(1696)* 4598GAT(1719)* ; 4654GAT(1745)
g1715 and 4531GAT(1698)* 4595GAT(1720)* ; 4650GAT(1746)
g1716 and 4526GAT(1700)* 4592GAT(1721)* ; 4646GAT(1747)
g1717 and 4704GAT(1725)* 1299GAT(35)* ; 4758GAT(1748)
g1718 and 4643GAT(1702)* 4704GAT(1725)* ; 4759GAT(1749)
g1719 and 4698GAT(1727)* 4701GAT(1726)* ; 4754GAT(1750)
g1720 and 4697GAT(1738)* 4696GAT(1728)* ; 4751GAT(1751)
g1721 and 4692GAT(1739)* 4515GAT(1649)* ; 4748GAT(1752)
g1722 and 4692GAT(1739)* 4634GAT(1704)* ; 4746GAT(1753)
g1723 and 4688GAT(1731)* 4687GAT(1730)* ; 4739GAT(1754)
g1724 and 4683GAT(1732)* 4625GAT(1708)* ; 4737GAT(1755)
g1725 and 4622GAT(1709)* 4683GAT(1732)* ; 4738GAT(1756)
g1726 and 4677GAT(1734)* 4680GAT(1733)* ; 4733GAT(1757)
g1727 and 4676GAT(1740)* 4675GAT(1735)* ; 4730GAT(1758)
g1728 and 4671GAT(1741)* 4494GAT(1656)* ; 4727GAT(1759)
g1729 and 4671GAT(1741)* 4613GAT(1711)* ; 4725GAT(1760)
g1730 and 4667GAT(1742)* 4666GAT(1737)* ; 4718GAT(1761)
g1731 and 4662GAT(1743)* 4604GAT(1715)* ; 4716GAT(1762)
g1732 and 4658GAT(1744)* 4601GAT(1717)* ; 4714GAT(1763)
g1733 and 4654GAT(1745)* 4598GAT(1719)* ; 4712GAT(1764)
g1734 and 1155GAT(83)* 4692GAT(1739)* ; 4747GAT(1765)
g1735 and 4650GAT(1746)* 4595GAT(1720)* ; 4710GAT(1766)
g1736 and 1107GAT(99)* 4689GAT(1729)* ; 4742GAT(1767)
g1737 and 4646GAT(1747)* 4592GAT(1721)* ; 4708GAT(1768)
g1738 and 912GAT(164)* 4671GAT(1741)* ; 4726GAT(1769)
g1739 and 864GAT(180)* 4668GAT(1736)* ; 4721GAT(1770)
g1740 and 4546GAT(1692)* 4662GAT(1743)* ; 4717GAT(1771)
g1741 and 4541GAT(1694)* 4658GAT(1744)* ; 4715GAT(1772)
g1742 and 4536GAT(1696)* 4654GAT(1745)* ; 4713GAT(1773)
g1743 and 4531GAT(1698)* 4650GAT(1746)* ; 4711GAT(1774)
g1744 and 4526GAT(1700)* 4646GAT(1747)* ; 4709GAT(1775)
g1745 and 4759GAT(1749)* 4758GAT(1748)* ; 4814GAT(1776)
g1746 and 4754GAT(1750)* 4701GAT(1726)* ; 4812GAT(1777)
g1747 and 4698GAT(1727)* 4754GAT(1750)* ; 4813GAT(1778)
g1748 and 4748GAT(1752)* 4751GAT(1751)* ; 4808GAT(1779)
g1749 and 4747GAT(1765)* 4746GAT(1753)* ; 4805GAT(1780)
g1750 and 4742GAT(1767)* 4578GAT(1672)* ; 4802GAT(1781)
g1751 and 4742GAT(1767)* 4689GAT(1729)* ; 4800GAT(1782)
g1752 and 4738GAT(1756)* 4737GAT(1755)* ; 4793GAT(1783)
g1753 and 4733GAT(1757)* 4680GAT(1733)* ; 4791GAT(1784)
g1754 and 4677GAT(1734)* 4733GAT(1757)* ; 4792GAT(1785)
g1755 and 4727GAT(1759)* 4730GAT(1758)* ; 4787GAT(1786)
g1756 and 4726GAT(1769)* 4725GAT(1760)* ; 4784GAT(1787)
g1757 and 4721GAT(1770)* 4557GAT(1679)* ; 4781GAT(1788)
g1758 and 4721GAT(1770)* 4668GAT(1736)* ; 4779GAT(1789)
g1759 and 4717GAT(1771)* 4716GAT(1762)* ; 4772GAT(1790)
g1760 and 4715GAT(1772)* 4714GAT(1763)* ; 4769GAT(1791)
g1761 and 4713GAT(1773)* 4712GAT(1764)* ; 4766GAT(1792)
g1762 and 4711GAT(1774)* 4710GAT(1766)* ; 4763GAT(1793)
g1763 and 1107GAT(99)* 4742GAT(1767)* ; 4801GAT(1794)
g1764 and 4709GAT(1775)* 4708GAT(1768)* ; 4760GAT(1795)
g1765 and 1059GAT(115)* 4739GAT(1754)* ; 4796GAT(1796)
g1766 and 864GAT(180)* 4721GAT(1770)* ; 4780GAT(1797)
g1767 and 816GAT(196)* 4718GAT(1761)* ; 4775GAT(1798)
g1768 and 4813GAT(1778)* 4812GAT(1777)* ; 4872GAT(1799)
g1769 and 4808GAT(1779)* 4751GAT(1751)* ; 4870GAT(1800)
g1770 and 4748GAT(1752)* 4808GAT(1779)* ; 4871GAT(1801)
g1771 and 4802GAT(1781)* 4805GAT(1780)* ; 4866GAT(1802)
g1772 and 4801GAT(1794)* 4800GAT(1782)* ; 4863GAT(1803)
g1773 and 4796GAT(1796)* 4628GAT(1707)* ; 4860GAT(1804)
g1774 and 4796GAT(1796)* 4739GAT(1754)* ; 4858GAT(1805)
g1775 and 4792GAT(1785)* 4791GAT(1784)* ; 4851GAT(1806)
g1776 and 4787GAT(1786)* 4730GAT(1758)* ; 4849GAT(1807)
g1777 and 4727GAT(1759)* 4787GAT(1786)* ; 4850GAT(1808)
g1778 and 4781GAT(1788)* 4784GAT(1787)* ; 4845GAT(1809)
g1779 and 4780GAT(1797)* 4779GAT(1789)* ; 4842GAT(1810)
g1780 and 4775GAT(1798)* 4607GAT(1714)* ; 4839GAT(1811)
g1781 and 4775GAT(1798)* 4718GAT(1761)* ; 4837GAT(1812)
g1782 and 1254GAT(50)* 4814GAT(1776)* ; 4875GAT(1813)
g1783 and 1059GAT(115)* 4796GAT(1796)* ; 4859GAT(1814)
g1784 and 1011GAT(131)* 4793GAT(1783)* ; 4854GAT(1815)
g1785 and 816GAT(196)* 4775GAT(1798)* ; 4838GAT(1816)
g1786 and 768GAT(212)* 4772GAT(1790)* ; 4833GAT(1817)
g1787 and 720GAT(228)* 4769GAT(1791)* ; 4829GAT(1818)
g1788 and 672GAT(244)* 4766GAT(1792)* ; 4825GAT(1819)
g1789 and 624GAT(260)* 4763GAT(1793)* ; 4821GAT(1820)
g1790 and 576GAT(276)* 4760GAT(1795)* ; 4817GAT(1821)
g1791 and 4875GAT(1813)* 4704GAT(1725)* ; 4943GAT(1822)
g1792 and 4875GAT(1813)* 4814GAT(1776)* ; 4941GAT(1823)
g1793 and 4871GAT(1801)* 4870GAT(1800)* ; 4934GAT(1824)
g1794 and 4866GAT(1802)* 4805GAT(1780)* ; 4932GAT(1825)
g1795 and 4802GAT(1781)* 4866GAT(1802)* ; 4933GAT(1826)
g1796 and 4860GAT(1804)* 4863GAT(1803)* ; 4928GAT(1827)
g1797 and 4859GAT(1814)* 4858GAT(1805)* ; 4925GAT(1828)
g1798 and 4854GAT(1815)* 4683GAT(1732)* ; 4922GAT(1829)
g1799 and 4854GAT(1815)* 4793GAT(1783)* ; 4920GAT(1830)
g1800 and 4850GAT(1808)* 4849GAT(1807)* ; 4913GAT(1831)
g1801 and 4845GAT(1809)* 4784GAT(1787)* ; 4911GAT(1832)
g1802 and 4781GAT(1788)* 4845GAT(1809)* ; 4912GAT(1833)
g1803 and 4839GAT(1811)* 4842GAT(1810)* ; 4907GAT(1834)
g1804 and 4838GAT(1816)* 4837GAT(1812)* ; 4904GAT(1835)
g1805 and 4833GAT(1817)* 4772GAT(1790)* ; 4899GAT(1836)
g1806 and 1254GAT(50)* 4875GAT(1813)* ; 4942GAT(1837)
g1807 and 4829GAT(1818)* 4769GAT(1791)* ; 4894GAT(1838)
g1808 and 1206GAT(66)* 4872GAT(1799)* ; 4937GAT(1839)
g1809 and 4825GAT(1819)* 4766GAT(1792)* ; 4889GAT(1840)
g1810 and 4821GAT(1820)* 4763GAT(1793)* ; 4884GAT(1841)
g1811 and 4817GAT(1821)* 4760GAT(1795)* ; 4879GAT(1842)
g1812 and 1011GAT(131)* 4854GAT(1815)* ; 4921GAT(1843)
g1813 and 963GAT(147)* 4851GAT(1806)* ; 4916GAT(1844)
g1814 and 4833GAT(1817)* 4662GAT(1743)* ; 4901GAT(1845)
g1815 and 768GAT(212)* 4833GAT(1817)* ; 4900GAT(1846)
g1816 and 4829GAT(1818)* 4658GAT(1744)* ; 4896GAT(1847)
g1817 and 720GAT(228)* 4829GAT(1818)* ; 4895GAT(1848)
g1818 and 4825GAT(1819)* 4654GAT(1745)* ; 4891GAT(1849)
g1819 and 672GAT(244)* 4825GAT(1819)* ; 4890GAT(1850)
g1820 and 4821GAT(1820)* 4650GAT(1746)* ; 4886GAT(1851)
g1821 and 624GAT(260)* 4821GAT(1820)* ; 4885GAT(1852)
g1822 and 4817GAT(1821)* 4646GAT(1747)* ; 4881GAT(1853)
g1823 and 576GAT(276)* 4817GAT(1821)* ; 4880GAT(1854)
g1824 and 4943GAT(1822)* 1302GAT(34)* ; 5001GAT(1855)
g1825 and 4942GAT(1837)* 4941GAT(1823)* ; 4998GAT(1856)
g1826 and 4937GAT(1839)* 4754GAT(1750)* ; 4995GAT(1857)
g1827 and 4937GAT(1839)* 4872GAT(1799)* ; 4993GAT(1858)
g1828 and 4933GAT(1826)* 4932GAT(1825)* ; 4986GAT(1859)
g1829 and 4928GAT(1827)* 4863GAT(1803)* ; 4984GAT(1860)
g1830 and 4860GAT(1804)* 4928GAT(1827)* ; 4985GAT(1861)
g1831 and 4922GAT(1829)* 4925GAT(1828)* ; 4980GAT(1862)
g1832 and 4921GAT(1843)* 4920GAT(1830)* ; 4977GAT(1863)
g1833 and 4916GAT(1844)* 4733GAT(1757)* ; 4974GAT(1864)
g1834 and 4916GAT(1844)* 4851GAT(1806)* ; 4972GAT(1865)
g1835 and 4912GAT(1833)* 4911GAT(1832)* ; 4965GAT(1866)
g1836 and 4907GAT(1834)* 4842GAT(1810)* ; 4963GAT(1867)
g1837 and 4839GAT(1811)* 4907GAT(1834)* ; 4964GAT(1868)
g1838 and 4901GAT(1845)* 4904GAT(1835)* ; 4959GAT(1869)
g1839 and 4900GAT(1846)* 4899GAT(1836)* ; 4956GAT(1870)
g1840 and 4895GAT(1848)* 4894GAT(1838)* ; 4953GAT(1871)
g1841 and 1206GAT(66)* 4937GAT(1839)* ; 4994GAT(1872)
g1842 and 4890GAT(1850)* 4889GAT(1840)* ; 4950GAT(1873)
g1843 and 1158GAT(82)* 4934GAT(1824)* ; 4989GAT(1874)
g1844 and 4885GAT(1852)* 4884GAT(1841)* ; 4947GAT(1875)
g1845 and 4880GAT(1854)* 4879GAT(1842)* ; 4946GAT(1876)
g1846 and 963GAT(147)* 4916GAT(1844)* ; 4973GAT(1877)
g1847 and 915GAT(163)* 4913GAT(1831)* ; 4968GAT(1878)
g1848 and 5001GAT(1855)* 1302GAT(34)* ; 5063GAT(1879)
g1849 and 4943GAT(1822)* 5001GAT(1855)* ; 5064GAT(1880)
g1850 and 4995GAT(1857)* 4998GAT(1856)* ; 5059GAT(1881)
g1851 and 4994GAT(1872)* 4993GAT(1858)* ; 5056GAT(1882)
g1852 and 4989GAT(1874)* 4808GAT(1779)* ; 5053GAT(1883)
g1853 and 4989GAT(1874)* 4934GAT(1824)* ; 5051GAT(1884)
g1854 and 4985GAT(1861)* 4984GAT(1860)* ; 5044GAT(1885)
g1855 and 4980GAT(1862)* 4925GAT(1828)* ; 5042GAT(1886)
g1856 and 4922GAT(1829)* 4980GAT(1862)* ; 5043GAT(1887)
g1857 and 4974GAT(1864)* 4977GAT(1863)* ; 5038GAT(1888)
g1858 and 4973GAT(1877)* 4972GAT(1865)* ; 5035GAT(1889)
g1859 and 4968GAT(1878)* 4787GAT(1786)* ; 5032GAT(1890)
g1860 and 4968GAT(1878)* 4913GAT(1831)* ; 5030GAT(1891)
g1861 and 4964GAT(1868)* 4963GAT(1867)* ; 5023GAT(1892)
g1862 and 4959GAT(1869)* 4904GAT(1835)* ; 5021GAT(1893)
g1863 and 1158GAT(82)* 4989GAT(1874)* ; 5052GAT(1894)
g1864 and 1110GAT(98)* 4986GAT(1859)* ; 5047GAT(1895)
g1865 and 915GAT(163)* 4968GAT(1878)* ; 5031GAT(1896)
g1866 and 867GAT(179)* 4965GAT(1866)* ; 5026GAT(1897)
g1867 and 4901GAT(1845)* 4959GAT(1869)* ; 5022GAT(1898)
g1868 and 4896GAT(1847)* 4956GAT(1870)* ; 5017GAT(1899)
g1869 and 4891GAT(1849)* 4953GAT(1871)* ; 5013GAT(1900)
g1870 and 4886GAT(1851)* 4950GAT(1873)* ; 5009GAT(1901)
g1871 and 4881GAT(1853)* 4947GAT(1875)* ; 5005GAT(1902)
g1872 and 5064GAT(1880)* 5063GAT(1879)* ; 5115GAT(1903)
g1873 and 5059GAT(1881)* 4998GAT(1856)* ; 5113GAT(1904)
g1874 and 4995GAT(1857)* 5059GAT(1881)* ; 5114GAT(1905)
g1875 and 5053GAT(1883)* 5056GAT(1882)* ; 5109GAT(1906)
g1876 and 5052GAT(1894)* 5051GAT(1884)* ; 5106GAT(1907)
g1877 and 5047GAT(1895)* 4866GAT(1802)* ; 5103GAT(1908)
g1878 and 5047GAT(1895)* 4986GAT(1859)* ; 5101GAT(1909)
g1879 and 5043GAT(1887)* 5042GAT(1886)* ; 5094GAT(1910)
g1880 and 5038GAT(1888)* 4977GAT(1863)* ; 5092GAT(1911)
g1881 and 4974GAT(1864)* 5038GAT(1888)* ; 5093GAT(1912)
g1882 and 5032GAT(1890)* 5035GAT(1889)* ; 5088GAT(1913)
g1883 and 5031GAT(1896)* 5030GAT(1891)* ; 5085GAT(1914)
g1884 and 5026GAT(1897)* 4845GAT(1809)* ; 5082GAT(1915)
g1885 and 5026GAT(1897)* 4965GAT(1866)* ; 5080GAT(1916)
g1886 and 5022GAT(1898)* 5021GAT(1893)* ; 5073GAT(1917)
g1887 and 5017GAT(1899)* 4956GAT(1870)* ; 5071GAT(1918)
g1888 and 5013GAT(1900)* 4953GAT(1871)* ; 5069GAT(1919)
g1889 and 5009GAT(1901)* 4950GAT(1873)* ; 5067GAT(1920)
g1890 and 5005GAT(1902)* 4947GAT(1875)* ; 5065GAT(1921)
g1891 and 1110GAT(98)* 5047GAT(1895)* ; 5102GAT(1922)
g1892 and 1062GAT(114)* 5044GAT(1885)* ; 5097GAT(1923)
g1893 and 867GAT(179)* 5026GAT(1897)* ; 5081GAT(1924)
g1894 and 819GAT(195)* 5023GAT(1892)* ; 5076GAT(1925)
g1895 and 4896GAT(1847)* 5017GAT(1899)* ; 5072GAT(1926)
g1896 and 4891GAT(1849)* 5013GAT(1900)* ; 5070GAT(1927)
g1897 and 4886GAT(1851)* 5009GAT(1901)* ; 5068GAT(1928)
g1898 and 4881GAT(1853)* 5005GAT(1902)* ; 5066GAT(1929)
g1899 and 5114GAT(1905)* 5113GAT(1904)* ; 5169GAT(1930)
g1900 and 5109GAT(1906)* 5056GAT(1882)* ; 5167GAT(1931)
g1901 and 5053GAT(1883)* 5109GAT(1906)* ; 5168GAT(1932)
g1902 and 5103GAT(1908)* 5106GAT(1907)* ; 5163GAT(1933)
g1903 and 5102GAT(1922)* 5101GAT(1909)* ; 5160GAT(1934)
g1904 and 5097GAT(1923)* 4928GAT(1827)* ; 5157GAT(1935)
g1905 and 5097GAT(1923)* 5044GAT(1885)* ; 5155GAT(1936)
g1906 and 5093GAT(1912)* 5092GAT(1911)* ; 5148GAT(1937)
g1907 and 5088GAT(1913)* 5035GAT(1889)* ; 5146GAT(1938)
g1908 and 5032GAT(1890)* 5088GAT(1913)* ; 5147GAT(1939)
g1909 and 5082GAT(1915)* 5085GAT(1914)* ; 5142GAT(1940)
g1910 and 5081GAT(1924)* 5080GAT(1916)* ; 5139GAT(1941)
g1911 and 5076GAT(1925)* 4907GAT(1834)* ; 5136GAT(1942)
g1912 and 5076GAT(1925)* 5023GAT(1892)* ; 5134GAT(1943)
g1913 and 5072GAT(1926)* 5071GAT(1918)* ; 5127GAT(1944)
g1914 and 1257GAT(49)* 5115GAT(1903)* ; 5172GAT(1945)
g1915 and 5070GAT(1927)* 5069GAT(1919)* ; 5124GAT(1946)
g1916 and 5068GAT(1928)* 5067GAT(1920)* ; 5121GAT(1947)
g1917 and 5066GAT(1929)* 5065GAT(1921)* ; 5118GAT(1948)
g1918 and 1062GAT(114)* 5097GAT(1923)* ; 5156GAT(1949)
g1919 and 1014GAT(130)* 5094GAT(1910)* ; 5151GAT(1950)
g1920 and 819GAT(195)* 5076GAT(1925)* ; 5135GAT(1951)
g1921 and 771GAT(211)* 5073GAT(1917)* ; 5130GAT(1952)
g1922 and 5172GAT(1945)* 5001GAT(1855)* ; 5236GAT(1953)
g1923 and 5172GAT(1945)* 5115GAT(1903)* ; 5234GAT(1954)
g1924 and 5168GAT(1932)* 5167GAT(1931)* ; 5227GAT(1955)
g1925 and 5163GAT(1933)* 5106GAT(1907)* ; 5225GAT(1956)
g1926 and 5103GAT(1908)* 5163GAT(1933)* ; 5226GAT(1957)
g1927 and 5157GAT(1935)* 5160GAT(1934)* ; 5221GAT(1958)
g1928 and 5156GAT(1949)* 5155GAT(1936)* ; 5218GAT(1959)
g1929 and 5151GAT(1950)* 4980GAT(1862)* ; 5215GAT(1960)
g1930 and 5151GAT(1950)* 5094GAT(1910)* ; 5213GAT(1961)
g1931 and 5147GAT(1939)* 5146GAT(1938)* ; 5206GAT(1962)
g1932 and 5142GAT(1940)* 5085GAT(1914)* ; 5204GAT(1963)
g1933 and 5082GAT(1915)* 5142GAT(1940)* ; 5205GAT(1964)
g1934 and 5136GAT(1942)* 5139GAT(1941)* ; 5200GAT(1965)
g1935 and 5135GAT(1951)* 5134GAT(1943)* ; 5197GAT(1966)
g1936 and 5130GAT(1952)* 4959GAT(1869)* ; 5194GAT(1967)
g1937 and 5130GAT(1952)* 5073GAT(1917)* ; 5192GAT(1968)
g1938 and 1257GAT(49)* 5172GAT(1945)* ; 5235GAT(1969)
g1939 and 1209GAT(65)* 5169GAT(1930)* ; 5230GAT(1970)
g1940 and 1014GAT(130)* 5151GAT(1950)* ; 5214GAT(1971)
g1941 and 966GAT(146)* 5148GAT(1937)* ; 5209GAT(1972)
g1942 and 771GAT(211)* 5130GAT(1952)* ; 5193GAT(1973)
g1943 and 723GAT(227)* 5127GAT(1944)* ; 5188GAT(1974)
g1944 and 675GAT(243)* 5124GAT(1946)* ; 5184GAT(1975)
g1945 and 627GAT(259)* 5121GAT(1947)* ; 5180GAT(1976)
g1946 and 579GAT(275)* 5118GAT(1948)* ; 5176GAT(1977)
g1947 and 5236GAT(1953)* 1305GAT(33)* ; 5304GAT(1978)
g1948 and 5235GAT(1969)* 5234GAT(1954)* ; 5301GAT(1979)
g1949 and 5230GAT(1970)* 5059GAT(1881)* ; 5298GAT(1980)
g1950 and 5230GAT(1970)* 5169GAT(1930)* ; 5296GAT(1981)
g1951 and 5226GAT(1957)* 5225GAT(1956)* ; 5289GAT(1982)
g1952 and 5221GAT(1958)* 5160GAT(1934)* ; 5287GAT(1983)
g1953 and 5157GAT(1935)* 5221GAT(1958)* ; 5288GAT(1984)
g1954 and 5215GAT(1960)* 5218GAT(1959)* ; 5283GAT(1985)
g1955 and 5214GAT(1971)* 5213GAT(1961)* ; 5280GAT(1986)
g1956 and 5209GAT(1972)* 5038GAT(1888)* ; 5277GAT(1987)
g1957 and 5209GAT(1972)* 5148GAT(1937)* ; 5275GAT(1988)
g1958 and 5205GAT(1964)* 5204GAT(1963)* ; 5268GAT(1989)
g1959 and 5200GAT(1965)* 5139GAT(1941)* ; 5266GAT(1990)
g1960 and 5136GAT(1942)* 5200GAT(1965)* ; 5267GAT(1991)
g1961 and 5194GAT(1967)* 5197GAT(1966)* ; 5262GAT(1992)
g1962 and 5193GAT(1973)* 5192GAT(1968)* ; 5259GAT(1993)
g1963 and 5188GAT(1974)* 5127GAT(1944)* ; 5254GAT(1994)
g1964 and 5184GAT(1975)* 5124GAT(1946)* ; 5249GAT(1995)
g1965 and 1209GAT(65)* 5230GAT(1970)* ; 5297GAT(1996)
g1966 and 5180GAT(1976)* 5121GAT(1947)* ; 5244GAT(1997)
g1967 and 1161GAT(81)* 5227GAT(1955)* ; 5292GAT(1998)
g1968 and 5176GAT(1977)* 5118GAT(1948)* ; 5239GAT(1999)
g1969 and 966GAT(146)* 5209GAT(1972)* ; 5276GAT(2000)
g1970 and 918GAT(162)* 5206GAT(1962)* ; 5271GAT(2001)
g1971 and 5188GAT(1974)* 5017GAT(1899)* ; 5256GAT(2002)
g1972 and 723GAT(227)* 5188GAT(1974)* ; 5255GAT(2003)
g1973 and 5184GAT(1975)* 5013GAT(1900)* ; 5251GAT(2004)
g1974 and 675GAT(243)* 5184GAT(1975)* ; 5250GAT(2005)
g1975 and 5180GAT(1976)* 5009GAT(1901)* ; 5246GAT(2006)
g1976 and 627GAT(259)* 5180GAT(1976)* ; 5245GAT(2007)
g1977 and 5176GAT(1977)* 5005GAT(1902)* ; 5241GAT(2008)
g1978 and 579GAT(275)* 5176GAT(1977)* ; 5240GAT(2009)
g1979 and 5304GAT(1978)* 1305GAT(33)* ; 5364GAT(2010)
g1980 and 5236GAT(1953)* 5304GAT(1978)* ; 5365GAT(2011)
g1981 and 5298GAT(1980)* 5301GAT(1979)* ; 5360GAT(2012)
g1982 and 5297GAT(1996)* 5296GAT(1981)* ; 5357GAT(2013)
g1983 and 5292GAT(1998)* 5109GAT(1906)* ; 5354GAT(2014)
g1984 and 5292GAT(1998)* 5227GAT(1955)* ; 5352GAT(2015)
g1985 and 5288GAT(1984)* 5287GAT(1983)* ; 5345GAT(2016)
g1986 and 5283GAT(1985)* 5218GAT(1959)* ; 5343GAT(2017)
g1987 and 5215GAT(1960)* 5283GAT(1985)* ; 5344GAT(2018)
g1988 and 5277GAT(1987)* 5280GAT(1986)* ; 5339GAT(2019)
g1989 and 5276GAT(2000)* 5275GAT(1988)* ; 5336GAT(2020)
g1990 and 5271GAT(2001)* 5088GAT(1913)* ; 5333GAT(2021)
g1991 and 5271GAT(2001)* 5206GAT(1962)* ; 5331GAT(2022)
g1992 and 5267GAT(1991)* 5266GAT(1990)* ; 5324GAT(2023)
g1993 and 5262GAT(1992)* 5197GAT(1966)* ; 5322GAT(2024)
g1994 and 5194GAT(1967)* 5262GAT(1992)* ; 5323GAT(2025)
g1995 and 5256GAT(2002)* 5259GAT(1993)* ; 5318GAT(2026)
g1996 and 5255GAT(2003)* 5254GAT(1994)* ; 5315GAT(2027)
g1997 and 5250GAT(2005)* 5249GAT(1995)* ; 5312GAT(2028)
g1998 and 5245GAT(2007)* 5244GAT(1997)* ; 5309GAT(2029)
g1999 and 1161GAT(81)* 5292GAT(1998)* ; 5353GAT(2030)
g2000 and 5240GAT(2009)* 5239GAT(1999)* ; 5308GAT(2031)
g2001 and 1113GAT(97)* 5289GAT(1982)* ; 5348GAT(2032)
g2002 and 918GAT(162)* 5271GAT(2001)* ; 5332GAT(2033)
g2003 and 870GAT(178)* 5268GAT(1989)* ; 5327GAT(2034)
g2004 and 5365GAT(2011)* 5364GAT(2010)* ; 5422GAT(2035)
g2005 and 5360GAT(2012)* 5301GAT(1979)* ; 5420GAT(2036)
g2006 and 5298GAT(1980)* 5360GAT(2012)* ; 5421GAT(2037)
g2007 and 5354GAT(2014)* 5357GAT(2013)* ; 5416GAT(2038)
g2008 and 5353GAT(2030)* 5352GAT(2015)* ; 5413GAT(2039)
g2009 and 5348GAT(2032)* 5163GAT(1933)* ; 5410GAT(2040)
g2010 and 5348GAT(2032)* 5289GAT(1982)* ; 5408GAT(2041)
g2011 and 5344GAT(2018)* 5343GAT(2017)* ; 5401GAT(2042)
g2012 and 5339GAT(2019)* 5280GAT(1986)* ; 5399GAT(2043)
g2013 and 5277GAT(1987)* 5339GAT(2019)* ; 5400GAT(2044)
g2014 and 5333GAT(2021)* 5336GAT(2020)* ; 5395GAT(2045)
g2015 and 5332GAT(2033)* 5331GAT(2022)* ; 5392GAT(2046)
g2016 and 5327GAT(2034)* 5142GAT(1940)* ; 5389GAT(2047)
g2017 and 5327GAT(2034)* 5268GAT(1989)* ; 5387GAT(2048)
g2018 and 5323GAT(2025)* 5322GAT(2024)* ; 5380GAT(2049)
g2019 and 5318GAT(2026)* 5259GAT(1993)* ; 5378GAT(2050)
g2020 and 1113GAT(97)* 5348GAT(2032)* ; 5409GAT(2051)
g2021 and 1065GAT(113)* 5345GAT(2016)* ; 5404GAT(2052)
g2022 and 870GAT(178)* 5327GAT(2034)* ; 5388GAT(2053)
g2023 and 822GAT(194)* 5324GAT(2023)* ; 5383GAT(2054)
g2024 and 5256GAT(2002)* 5318GAT(2026)* ; 5379GAT(2055)
g2025 and 5251GAT(2004)* 5315GAT(2027)* ; 5374GAT(2056)
g2026 and 5246GAT(2006)* 5312GAT(2028)* ; 5370GAT(2057)
g2027 and 5241GAT(2008)* 5309GAT(2029)* ; 5366GAT(2058)
g2028 and 5421GAT(2037)* 5420GAT(2036)* ; 5473GAT(2059)
g2029 and 5416GAT(2038)* 5357GAT(2013)* ; 5471GAT(2060)
g2030 and 5354GAT(2014)* 5416GAT(2038)* ; 5472GAT(2061)
g2031 and 5410GAT(2040)* 5413GAT(2039)* ; 5467GAT(2062)
g2032 and 5409GAT(2051)* 5408GAT(2041)* ; 5464GAT(2063)
g2033 and 5404GAT(2052)* 5221GAT(1958)* ; 5461GAT(2064)
g2034 and 5404GAT(2052)* 5345GAT(2016)* ; 5459GAT(2065)
g2035 and 5400GAT(2044)* 5399GAT(2043)* ; 5452GAT(2066)
g2036 and 5395GAT(2045)* 5336GAT(2020)* ; 5450GAT(2067)
g2037 and 5333GAT(2021)* 5395GAT(2045)* ; 5451GAT(2068)
g2038 and 5389GAT(2047)* 5392GAT(2046)* ; 5446GAT(2069)
g2039 and 5388GAT(2053)* 5387GAT(2048)* ; 5443GAT(2070)
g2040 and 5383GAT(2054)* 5200GAT(1965)* ; 5440GAT(2071)
g2041 and 5383GAT(2054)* 5324GAT(2023)* ; 5438GAT(2072)
g2042 and 5379GAT(2055)* 5378GAT(2050)* ; 5431GAT(2073)
g2043 and 5374GAT(2056)* 5315GAT(2027)* ; 5429GAT(2074)
g2044 and 1260GAT(48)* 5422GAT(2035)* ; 5476GAT(2075)
g2045 and 5370GAT(2057)* 5312GAT(2028)* ; 5427GAT(2076)
g2046 and 5366GAT(2058)* 5309GAT(2029)* ; 5425GAT(2077)
g2047 and 1065GAT(113)* 5404GAT(2052)* ; 5460GAT(2078)
g2048 and 1017GAT(129)* 5401GAT(2042)* ; 5455GAT(2079)
g2049 and 822GAT(194)* 5383GAT(2054)* ; 5439GAT(2080)
g2050 and 774GAT(210)* 5380GAT(2049)* ; 5434GAT(2081)
g2051 and 5251GAT(2004)* 5374GAT(2056)* ; 5430GAT(2082)
g2052 and 5246GAT(2006)* 5370GAT(2057)* ; 5428GAT(2083)
g2053 and 5241GAT(2008)* 5366GAT(2058)* ; 5426GAT(2084)
g2054 and 5476GAT(2075)* 5304GAT(1978)* ; 5537GAT(2085)
g2055 and 5476GAT(2075)* 5422GAT(2035)* ; 5535GAT(2086)
g2056 and 5472GAT(2061)* 5471GAT(2060)* ; 5528GAT(2087)
g2057 and 5467GAT(2062)* 5413GAT(2039)* ; 5526GAT(2088)
g2058 and 5410GAT(2040)* 5467GAT(2062)* ; 5527GAT(2089)
g2059 and 5461GAT(2064)* 5464GAT(2063)* ; 5522GAT(2090)
g2060 and 5460GAT(2078)* 5459GAT(2065)* ; 5519GAT(2091)
g2061 and 5455GAT(2079)* 5283GAT(1985)* ; 5516GAT(2092)
g2062 and 5455GAT(2079)* 5401GAT(2042)* ; 5514GAT(2093)
g2063 and 5451GAT(2068)* 5450GAT(2067)* ; 5507GAT(2094)
g2064 and 5446GAT(2069)* 5392GAT(2046)* ; 5505GAT(2095)
g2065 and 5389GAT(2047)* 5446GAT(2069)* ; 5506GAT(2096)
g2066 and 5440GAT(2071)* 5443GAT(2070)* ; 5501GAT(2097)
g2067 and 5439GAT(2080)* 5438GAT(2072)* ; 5498GAT(2098)
g2068 and 5434GAT(2081)* 5262GAT(1992)* ; 5495GAT(2099)
g2069 and 5434GAT(2081)* 5380GAT(2049)* ; 5493GAT(2100)
g2070 and 5430GAT(2082)* 5429GAT(2074)* ; 5486GAT(2101)
g2071 and 1260GAT(48)* 5476GAT(2075)* ; 5536GAT(2102)
g2072 and 5428GAT(2083)* 5427GAT(2076)* ; 5483GAT(2103)
g2073 and 1212GAT(64)* 5473GAT(2059)* ; 5531GAT(2104)
g2074 and 5426GAT(2084)* 5425GAT(2077)* ; 5480GAT(2105)
g2075 and 1017GAT(129)* 5455GAT(2079)* ; 5515GAT(2106)
g2076 and 969GAT(145)* 5452GAT(2066)* ; 5510GAT(2107)
g2077 and 774GAT(210)* 5434GAT(2081)* ; 5494GAT(2108)
g2078 and 726GAT(226)* 5431GAT(2073)* ; 5489GAT(2109)
g2079 and 5537GAT(2085)* 1308GAT(32)* ; 5602GAT(2110)
g2080 and 5536GAT(2102)* 5535GAT(2086)* ; 5599GAT(2111)
g2081 and 5531GAT(2104)* 5360GAT(2012)* ; 5596GAT(2112)
g2082 and 5531GAT(2104)* 5473GAT(2059)* ; 5594GAT(2113)
g2083 and 5527GAT(2089)* 5526GAT(2088)* ; 5587GAT(2114)
g2084 and 5522GAT(2090)* 5464GAT(2063)* ; 5585GAT(2115)
g2085 and 5461GAT(2064)* 5522GAT(2090)* ; 5586GAT(2116)
g2086 and 5516GAT(2092)* 5519GAT(2091)* ; 5581GAT(2117)
g2087 and 5515GAT(2106)* 5514GAT(2093)* ; 5578GAT(2118)
g2088 and 5510GAT(2107)* 5339GAT(2019)* ; 5575GAT(2119)
g2089 and 5510GAT(2107)* 5452GAT(2066)* ; 5573GAT(2120)
g2090 and 5506GAT(2096)* 5505GAT(2095)* ; 5566GAT(2121)
g2091 and 5501GAT(2097)* 5443GAT(2070)* ; 5564GAT(2122)
g2092 and 5440GAT(2071)* 5501GAT(2097)* ; 5565GAT(2123)
g2093 and 5495GAT(2099)* 5498GAT(2098)* ; 5560GAT(2124)
g2094 and 5494GAT(2108)* 5493GAT(2100)* ; 5557GAT(2125)
g2095 and 5489GAT(2109)* 5318GAT(2026)* ; 5554GAT(2126)
g2096 and 5489GAT(2109)* 5431GAT(2073)* ; 5552GAT(2127)
g2097 and 1212GAT(64)* 5531GAT(2104)* ; 5595GAT(2128)
g2098 and 1164GAT(80)* 5528GAT(2087)* ; 5590GAT(2129)
g2099 and 969GAT(145)* 5510GAT(2107)* ; 5574GAT(2130)
g2100 and 921GAT(161)* 5507GAT(2094)* ; 5569GAT(2131)
g2101 and 726GAT(226)* 5489GAT(2109)* ; 5553GAT(2132)
g2102 and 678GAT(242)* 5486GAT(2101)* ; 5548GAT(2133)
g2103 and 630GAT(258)* 5483GAT(2103)* ; 5544GAT(2134)
g2104 and 582GAT(274)* 5480GAT(2105)* ; 5540GAT(2135)
g2105 and 5602GAT(2110)* 1308GAT(32)* ; 5670GAT(2136)
g2106 and 5537GAT(2085)* 5602GAT(2110)* ; 5671GAT(2137)
g2107 and 5596GAT(2112)* 5599GAT(2111)* ; 5666GAT(2138)
g2108 and 5595GAT(2128)* 5594GAT(2113)* ; 5663GAT(2139)
g2109 and 5590GAT(2129)* 5416GAT(2038)* ; 5660GAT(2140)
g2110 and 5590GAT(2129)* 5528GAT(2087)* ; 5658GAT(2141)
g2111 and 5586GAT(2116)* 5585GAT(2115)* ; 5651GAT(2142)
g2112 and 5581GAT(2117)* 5519GAT(2091)* ; 5649GAT(2143)
g2113 and 5516GAT(2092)* 5581GAT(2117)* ; 5650GAT(2144)
g2114 and 5575GAT(2119)* 5578GAT(2118)* ; 5645GAT(2145)
g2115 and 5574GAT(2130)* 5573GAT(2120)* ; 5642GAT(2146)
g2116 and 5569GAT(2131)* 5395GAT(2045)* ; 5639GAT(2147)
g2117 and 5569GAT(2131)* 5507GAT(2094)* ; 5637GAT(2148)
g2118 and 5565GAT(2123)* 5564GAT(2122)* ; 5630GAT(2149)
g2119 and 5560GAT(2124)* 5498GAT(2098)* ; 5628GAT(2150)
g2120 and 5495GAT(2099)* 5560GAT(2124)* ; 5629GAT(2151)
g2121 and 5554GAT(2126)* 5557GAT(2125)* ; 5624GAT(2152)
g2122 and 5553GAT(2132)* 5552GAT(2127)* ; 5621GAT(2153)
g2123 and 5548GAT(2133)* 5486GAT(2101)* ; 5616GAT(2154)
g2124 and 5544GAT(2134)* 5483GAT(2103)* ; 5611GAT(2155)
g2125 and 5540GAT(2135)* 5480GAT(2105)* ; 5606GAT(2156)
g2126 and 1164GAT(80)* 5590GAT(2129)* ; 5659GAT(2157)
g2127 and 1116GAT(96)* 5587GAT(2114)* ; 5654GAT(2158)
g2128 and 921GAT(161)* 5569GAT(2131)* ; 5638GAT(2159)
g2129 and 873GAT(177)* 5566GAT(2121)* ; 5633GAT(2160)
g2130 and 5548GAT(2133)* 5374GAT(2056)* ; 5618GAT(2161)
g2131 and 678GAT(242)* 5548GAT(2133)* ; 5617GAT(2162)
g2132 and 5544GAT(2134)* 5370GAT(2057)* ; 5613GAT(2163)
g2133 and 630GAT(258)* 5544GAT(2134)* ; 5612GAT(2164)
g2134 and 5540GAT(2135)* 5366GAT(2058)* ; 5608GAT(2165)
g2135 and 582GAT(274)* 5540GAT(2135)* ; 5607GAT(2166)
g2136 and 5671GAT(2137)* 5670GAT(2136)* ; 5727GAT(2167)
g2137 and 5666GAT(2138)* 5599GAT(2111)* ; 5725GAT(2168)
g2138 and 5596GAT(2112)* 5666GAT(2138)* ; 5726GAT(2169)
g2139 and 5660GAT(2140)* 5663GAT(2139)* ; 5721GAT(2170)
g2140 and 5659GAT(2157)* 5658GAT(2141)* ; 5718GAT(2171)
g2141 and 5654GAT(2158)* 5467GAT(2062)* ; 5715GAT(2172)
g2142 and 5654GAT(2158)* 5587GAT(2114)* ; 5713GAT(2173)
g2143 and 5650GAT(2144)* 5649GAT(2143)* ; 5706GAT(2174)
g2144 and 5645GAT(2145)* 5578GAT(2118)* ; 5704GAT(2175)
g2145 and 5575GAT(2119)* 5645GAT(2145)* ; 5705GAT(2176)
g2146 and 5639GAT(2147)* 5642GAT(2146)* ; 5700GAT(2177)
g2147 and 5638GAT(2159)* 5637GAT(2148)* ; 5697GAT(2178)
g2148 and 5633GAT(2160)* 5446GAT(2069)* ; 5694GAT(2179)
g2149 and 5633GAT(2160)* 5566GAT(2121)* ; 5692GAT(2180)
g2150 and 5629GAT(2151)* 5628GAT(2150)* ; 5685GAT(2181)
g2151 and 5624GAT(2152)* 5557GAT(2125)* ; 5683GAT(2182)
g2152 and 5554GAT(2126)* 5624GAT(2152)* ; 5684GAT(2183)
g2153 and 5618GAT(2161)* 5621GAT(2153)* ; 5679GAT(2184)
g2154 and 5617GAT(2162)* 5616GAT(2154)* ; 5676GAT(2185)
g2155 and 5612GAT(2164)* 5611GAT(2155)* ; 5673GAT(2186)
g2156 and 5607GAT(2166)* 5606GAT(2156)* ; 5672GAT(2187)
g2157 and 1116GAT(96)* 5654GAT(2158)* ; 5714GAT(2188)
g2158 and 1068GAT(112)* 5651GAT(2142)* ; 5709GAT(2189)
g2159 and 873GAT(177)* 5633GAT(2160)* ; 5693GAT(2190)
g2160 and 825GAT(193)* 5630GAT(2149)* ; 5688GAT(2191)
g2161 and 5726GAT(2169)* 5725GAT(2168)* ; 5782GAT(2192)
g2162 and 5721GAT(2170)* 5663GAT(2139)* ; 5780GAT(2193)
g2163 and 5660GAT(2140)* 5721GAT(2170)* ; 5781GAT(2194)
g2164 and 5715GAT(2172)* 5718GAT(2171)* ; 5776GAT(2195)
g2165 and 5714GAT(2188)* 5713GAT(2173)* ; 5773GAT(2196)
g2166 and 5709GAT(2189)* 5522GAT(2090)* ; 5770GAT(2197)
g2167 and 5709GAT(2189)* 5651GAT(2142)* ; 5768GAT(2198)
g2168 and 5705GAT(2176)* 5704GAT(2175)* ; 5761GAT(2199)
g2169 and 5700GAT(2177)* 5642GAT(2146)* ; 5759GAT(2200)
g2170 and 5639GAT(2147)* 5700GAT(2177)* ; 5760GAT(2201)
g2171 and 5694GAT(2179)* 5697GAT(2178)* ; 5755GAT(2202)
g2172 and 5693GAT(2190)* 5692GAT(2180)* ; 5752GAT(2203)
g2173 and 5688GAT(2191)* 5501GAT(2097)* ; 5749GAT(2204)
g2174 and 5688GAT(2191)* 5630GAT(2149)* ; 5747GAT(2205)
g2175 and 5684GAT(2183)* 5683GAT(2182)* ; 5740GAT(2206)
g2176 and 5679GAT(2184)* 5621GAT(2153)* ; 5738GAT(2207)
g2177 and 1068GAT(112)* 5709GAT(2189)* ; 5769GAT(2208)
g2178 and 1020GAT(128)* 5706GAT(2174)* ; 5764GAT(2209)
g2179 and 825GAT(193)* 5688GAT(2191)* ; 5748GAT(2210)
g2180 and 777GAT(209)* 5685GAT(2181)* ; 5743GAT(2211)
g2181 and 5618GAT(2161)* 5679GAT(2184)* ; 5739GAT(2212)
g2182 and 5613GAT(2163)* 5676GAT(2185)* ; 5734GAT(2213)
g2183 and 5608GAT(2165)* 5673GAT(2186)* ; 5730GAT(2214)
g2184 and 5781GAT(2194)* 5780GAT(2193)* ; 5831GAT(2215)
g2185 and 5776GAT(2195)* 5718GAT(2171)* ; 5829GAT(2216)
g2186 and 5715GAT(2172)* 5776GAT(2195)* ; 5830GAT(2217)
g2187 and 5770GAT(2197)* 5773GAT(2196)* ; 5825GAT(2218)
g2188 and 5769GAT(2208)* 5768GAT(2198)* ; 5822GAT(2219)
g2189 and 5764GAT(2209)* 5581GAT(2117)* ; 5819GAT(2220)
g2190 and 5764GAT(2209)* 5706GAT(2174)* ; 5817GAT(2221)
g2191 and 5760GAT(2201)* 5759GAT(2200)* ; 5810GAT(2222)
g2192 and 5755GAT(2202)* 5697GAT(2178)* ; 5808GAT(2223)
g2193 and 5694GAT(2179)* 5755GAT(2202)* ; 5809GAT(2224)
g2194 and 5749GAT(2204)* 5752GAT(2203)* ; 5804GAT(2225)
g2195 and 5748GAT(2210)* 5747GAT(2205)* ; 5801GAT(2226)
g2196 and 5743GAT(2211)* 5560GAT(2124)* ; 5798GAT(2227)
g2197 and 5743GAT(2211)* 5685GAT(2181)* ; 5796GAT(2228)
g2198 and 5739GAT(2212)* 5738GAT(2207)* ; 5789GAT(2229)
g2199 and 5734GAT(2213)* 5676GAT(2185)* ; 5787GAT(2230)
g2200 and 5730GAT(2214)* 5673GAT(2186)* ; 5785GAT(2231)
g2201 and 1020GAT(128)* 5764GAT(2209)* ; 5818GAT(2232)
g2202 and 972GAT(144)* 5761GAT(2199)* ; 5813GAT(2233)
g2203 and 777GAT(209)* 5743GAT(2211)* ; 5797GAT(2234)
g2204 and 729GAT(225)* 5740GAT(2206)* ; 5792GAT(2235)
g2205 and 5613GAT(2163)* 5734GAT(2213)* ; 5788GAT(2236)
g2206 and 5608GAT(2165)* 5730GAT(2214)* ; 5786GAT(2237)
g2207 and 5830GAT(2217)* 5829GAT(2216)* ; 5879GAT(2238)
g2208 and 5825GAT(2218)* 5773GAT(2196)* ; 5877GAT(2239)
g2209 and 5770GAT(2197)* 5825GAT(2218)* ; 5878GAT(2240)
g2210 and 5819GAT(2220)* 5822GAT(2219)* ; 5873GAT(2241)
g2211 and 5818GAT(2232)* 5817GAT(2221)* ; 5870GAT(2242)
g2212 and 5813GAT(2233)* 5645GAT(2145)* ; 5867GAT(2243)
g2213 and 5813GAT(2233)* 5761GAT(2199)* ; 5865GAT(2244)
g2214 and 5809GAT(2224)* 5808GAT(2223)* ; 5858GAT(2245)
g2215 and 5804GAT(2225)* 5752GAT(2203)* ; 5856GAT(2246)
g2216 and 5749GAT(2204)* 5804GAT(2225)* ; 5857GAT(2247)
g2217 and 5798GAT(2227)* 5801GAT(2226)* ; 5852GAT(2248)
g2218 and 5797GAT(2234)* 5796GAT(2228)* ; 5849GAT(2249)
g2219 and 5792GAT(2235)* 5624GAT(2152)* ; 5846GAT(2250)
g2220 and 5792GAT(2235)* 5740GAT(2206)* ; 5844GAT(2251)
g2221 and 5788GAT(2236)* 5787GAT(2230)* ; 5837GAT(2252)
g2222 and 5786GAT(2237)* 5785GAT(2231)* ; 5834GAT(2253)
g2223 and 972GAT(144)* 5813GAT(2233)* ; 5866GAT(2254)
g2224 and 924GAT(160)* 5810GAT(2222)* ; 5861GAT(2255)
g2225 and 729GAT(225)* 5792GAT(2235)* ; 5845GAT(2256)
g2226 and 681GAT(241)* 5789GAT(2229)* ; 5840GAT(2257)
g2227 and 5878GAT(2240)* 5877GAT(2239)* ; 5925GAT(2258)
g2228 and 5873GAT(2241)* 5822GAT(2219)* ; 5923GAT(2259)
g2229 and 5819GAT(2220)* 5873GAT(2241)* ; 5924GAT(2260)
g2230 and 5867GAT(2243)* 5870GAT(2242)* ; 5919GAT(2261)
g2231 and 5866GAT(2254)* 5865GAT(2244)* ; 5916GAT(2262)
g2232 and 5861GAT(2255)* 5700GAT(2177)* ; 5913GAT(2263)
g2233 and 5861GAT(2255)* 5810GAT(2222)* ; 5911GAT(2264)
g2234 and 5857GAT(2247)* 5856GAT(2246)* ; 5904GAT(2265)
g2235 and 5852GAT(2248)* 5801GAT(2226)* ; 5902GAT(2266)
g2236 and 5798GAT(2227)* 5852GAT(2248)* ; 5903GAT(2267)
g2237 and 5846GAT(2250)* 5849GAT(2249)* ; 5898GAT(2268)
g2238 and 5845GAT(2256)* 5844GAT(2251)* ; 5895GAT(2269)
g2239 and 5840GAT(2257)* 5679GAT(2184)* ; 5892GAT(2270)
g2240 and 5840GAT(2257)* 5789GAT(2229)* ; 5890GAT(2271)
g2241 and 924GAT(160)* 5861GAT(2255)* ; 5912GAT(2272)
g2242 and 876GAT(176)* 5858GAT(2245)* ; 5907GAT(2273)
g2243 and 681GAT(241)* 5840GAT(2257)* ; 5891GAT(2274)
g2244 and 633GAT(257)* 5837GAT(2252)* ; 5886GAT(2275)
g2245 and 585GAT(273)* 5834GAT(2253)* ; 5882GAT(2276)
g2246 and 5924GAT(2260)* 5923GAT(2259)* ; 5968GAT(2277)
g2247 and 5919GAT(2261)* 5870GAT(2242)* ; 5966GAT(2278)
g2248 and 5867GAT(2243)* 5919GAT(2261)* ; 5967GAT(2279)
g2249 and 5913GAT(2263)* 5916GAT(2262)* ; 5962GAT(2280)
g2250 and 5912GAT(2272)* 5911GAT(2264)* ; 5959GAT(2281)
g2251 and 5907GAT(2273)* 5755GAT(2202)* ; 5956GAT(2282)
g2252 and 5907GAT(2273)* 5858GAT(2245)* ; 5954GAT(2283)
g2253 and 5903GAT(2267)* 5902GAT(2266)* ; 5947GAT(2284)
g2254 and 5898GAT(2268)* 5849GAT(2249)* ; 5945GAT(2285)
g2255 and 5846GAT(2250)* 5898GAT(2268)* ; 5946GAT(2286)
g2256 and 5892GAT(2270)* 5895GAT(2269)* ; 5941GAT(2287)
g2257 and 5891GAT(2274)* 5890GAT(2271)* ; 5938GAT(2288)
g2258 and 5886GAT(2275)* 5837GAT(2252)* ; 5933GAT(2289)
g2259 and 5882GAT(2276)* 5834GAT(2253)* ; 5928GAT(2290)
g2260 and 876GAT(176)* 5907GAT(2273)* ; 5955GAT(2291)
g2261 and 828GAT(192)* 5904GAT(2265)* ; 5950GAT(2292)
g2262 and 5886GAT(2275)* 5734GAT(2213)* ; 5935GAT(2293)
g2263 and 633GAT(257)* 5886GAT(2275)* ; 5934GAT(2294)
g2264 and 5882GAT(2276)* 5730GAT(2214)* ; 5930GAT(2295)
g2265 and 585GAT(273)* 5882GAT(2276)* ; 5929GAT(2296)
g2266 and 5967GAT(2279)* 5966GAT(2278)* ; 6002GAT(2297)
g2267 and 5962GAT(2280)* 5916GAT(2262)* ; 6000GAT(2298)
g2268 and 5913GAT(2263)* 5962GAT(2280)* ; 6001GAT(2299)
g2269 and 5956GAT(2282)* 5959GAT(2281)* ; 5996GAT(2300)
g2270 and 5955GAT(2291)* 5954GAT(2283)* ; 5993GAT(2301)
g2271 and 5950GAT(2292)* 5804GAT(2225)* ; 5990GAT(2302)
g2272 and 5950GAT(2292)* 5904GAT(2265)* ; 5988GAT(2303)
g2273 and 5946GAT(2286)* 5945GAT(2285)* ; 5981GAT(2304)
g2274 and 5941GAT(2287)* 5895GAT(2269)* ; 5979GAT(2305)
g2275 and 5892GAT(2270)* 5941GAT(2287)* ; 5980GAT(2306)
g2276 and 5935GAT(2293)* 5938GAT(2288)* ; 5975GAT(2307)
g2277 and 5934GAT(2294)* 5933GAT(2289)* ; 5972GAT(2308)
g2278 and 5929GAT(2296)* 5928GAT(2290)* ; 5971GAT(2309)
g2279 and 828GAT(192)* 5950GAT(2292)* ; 5989GAT(2310)
g2280 and 780GAT(208)* 5947GAT(2284)* ; 5984GAT(2311)
g2281 and 6001GAT(2299)* 6000GAT(2298)* ; 6032GAT(2312)
g2282 and 5996GAT(2300)* 5959GAT(2281)* ; 6030GAT(2313)
g2283 and 5956GAT(2282)* 5996GAT(2300)* ; 6031GAT(2314)
g2284 and 5990GAT(2302)* 5993GAT(2301)* ; 6026GAT(2315)
g2285 and 5989GAT(2310)* 5988GAT(2303)* ; 6023GAT(2316)
g2286 and 5984GAT(2311)* 5852GAT(2248)* ; 6020GAT(2317)
g2287 and 5984GAT(2311)* 5947GAT(2284)* ; 6018GAT(2318)
g2288 and 5980GAT(2306)* 5979GAT(2305)* ; 6011GAT(2319)
g2289 and 5975GAT(2307)* 5938GAT(2288)* ; 6009GAT(2320)
g2290 and 780GAT(208)* 5984GAT(2311)* ; 6019GAT(2321)
g2291 and 732GAT(224)* 5981GAT(2304)* ; 6014GAT(2322)
g2292 and 5935GAT(2293)* 5975GAT(2307)* ; 6010GAT(2323)
g2293 and 5930GAT(2295)* 5972GAT(2308)* ; 6005GAT(2324)
g2294 and 6031GAT(2314)* 6030GAT(2313)* ; 6058GAT(2325)
g2295 and 6026GAT(2315)* 5993GAT(2301)* ; 6056GAT(2326)
g2296 and 5990GAT(2302)* 6026GAT(2315)* ; 6057GAT(2327)
g2297 and 6020GAT(2317)* 6023GAT(2316)* ; 6052GAT(2328)
g2298 and 6019GAT(2321)* 6018GAT(2318)* ; 6049GAT(2329)
g2299 and 6014GAT(2322)* 5898GAT(2268)* ; 6046GAT(2330)
g2300 and 6014GAT(2322)* 5981GAT(2304)* ; 6044GAT(2331)
g2301 and 6010GAT(2323)* 6009GAT(2320)* ; 6037GAT(2332)
g2302 and 6005GAT(2324)* 5972GAT(2308)* ; 6035GAT(2333)
g2303 and 732GAT(224)* 6014GAT(2322)* ; 6045GAT(2334)
g2304 and 684GAT(240)* 6011GAT(2319)* ; 6040GAT(2335)
g2305 and 5930GAT(2295)* 6005GAT(2324)* ; 6036GAT(2336)
g2306 and 6057GAT(2327)* 6056GAT(2326)* ; 6082GAT(2337)
g2307 and 6052GAT(2328)* 6023GAT(2316)* ; 6080GAT(2338)
g2308 and 6020GAT(2317)* 6052GAT(2328)* ; 6081GAT(2339)
g2309 and 6046GAT(2330)* 6049GAT(2329)* ; 6076GAT(2340)
g2310 and 6045GAT(2334)* 6044GAT(2331)* ; 6073GAT(2341)
g2311 and 6040GAT(2335)* 5941GAT(2287)* ; 6070GAT(2342)
g2312 and 6040GAT(2335)* 6011GAT(2319)* ; 6068GAT(2343)
g2313 and 6036GAT(2336)* 6035GAT(2333)* ; 6061GAT(2344)
g2314 and 684GAT(240)* 6040GAT(2335)* ; 6069GAT(2345)
g2315 and 636GAT(256)* 6037GAT(2332)* ; 6064GAT(2346)
g2316 and 6081GAT(2339)* 6080GAT(2338)* ; 6103GAT(2347)
g2317 and 6076GAT(2340)* 6049GAT(2329)* ; 6101GAT(2348)
g2318 and 6046GAT(2330)* 6076GAT(2340)* ; 6102GAT(2349)
g2319 and 6070GAT(2342)* 6073GAT(2341)* ; 6097GAT(2350)
g2320 and 6069GAT(2345)* 6068GAT(2343)* ; 6094GAT(2351)
g2321 and 6064GAT(2346)* 5975GAT(2307)* ; 6091GAT(2352)
g2322 and 6064GAT(2346)* 6037GAT(2332)* ; 6089GAT(2353)
g2323 and 636GAT(256)* 6064GAT(2346)* ; 6090GAT(2354)
g2324 and 588GAT(272)* 6061GAT(2344)* ; 6085GAT(2355)
g2325 and 6102GAT(2349)* 6101GAT(2348)* ; 6120GAT(2356)
g2326 and 6097GAT(2350)* 6073GAT(2341)* ; 6118GAT(2357)
g2327 and 6070GAT(2342)* 6097GAT(2350)* ; 6119GAT(2358)
g2328 and 6091GAT(2352)* 6094GAT(2351)* ; 6114GAT(2359)
g2329 and 6090GAT(2354)* 6089GAT(2353)* ; 6111GAT(2360)
g2330 and 6085GAT(2355)* 6061GAT(2344)* ; 6106GAT(2361)
g2331 and 6085GAT(2355)* 6005GAT(2324)* ; 6108GAT(2362)
g2332 and 588GAT(272)* 6085GAT(2355)* ; 6107GAT(2363)
g2333 and 6119GAT(2358)* 6118GAT(2357)* ; 6130GAT(2364)
g2334 and 6114GAT(2359)* 6094GAT(2351)* ; 6128GAT(2365)
g2335 and 6091GAT(2352)* 6114GAT(2359)* ; 6129GAT(2366)
g2336 and 6108GAT(2362)* 6111GAT(2360)* ; 6124GAT(2367)
g2337 and 6107GAT(2363)* 6106GAT(2361)* ; 6123GAT(2368)
g2338 and 6129GAT(2366)* 6128GAT(2365)* ; 6135GAT(2369)
g2339 and 6124GAT(2367)* 6111GAT(2360)* ; 6133GAT(2370)
g2340 and 6108GAT(2362)* 6124GAT(2367)* ; 6134GAT(2371)
g2341 and 6134GAT(2371)* 6133GAT(2370)* ; 6138GAT(2372)
g2342 and 6138GAT(2372) ; 6141GAT(2373)
g2343 and 6141GAT(2373)* 6124GAT(2367)* ; 6147GAT(2374)
g2344 and 6141GAT(2373)* 6138GAT(2372)* ; 6145GAT(2375)
g2345 and 6141GAT(2373) ; 6146GAT(2376)
g2346 and 6147GAT(2374)* 6135GAT(2369)* ; 6151GAT(2377)
g2347 and 6146GAT(2376)* 6145GAT(2375)* ; 6150GAT(2378)
g2348 and 6151GAT(2377)* 6114GAT(2359)* ; 6157GAT(2379)
g2349 and 6151GAT(2377)* 6135GAT(2369)* ; 6155GAT(2380)
g2350 and 6147GAT(2374)* 6151GAT(2377)* ; 6156GAT(2381)
g2351 and 6157GAT(2379)* 6130GAT(2364)* ; 6161GAT(2382)
g2352 and 6156GAT(2381)* 6155GAT(2380)* ; 6160GAT(2383)
g2353 and 6161GAT(2382)* 6097GAT(2350)* ; 6167GAT(2384)
g2354 and 6161GAT(2382)* 6130GAT(2364)* ; 6165GAT(2385)
g2355 and 6157GAT(2379)* 6161GAT(2382)* ; 6166GAT(2386)
g2356 and 6167GAT(2384)* 6120GAT(2356)* ; 6171GAT(2387)
g2357 and 6166GAT(2386)* 6165GAT(2385)* ; 6170GAT(2388)
g2358 and 6171GAT(2387)* 6076GAT(2340)* ; 6177GAT(2389)
g2359 and 6171GAT(2387)* 6120GAT(2356)* ; 6175GAT(2390)
g2360 and 6167GAT(2384)* 6171GAT(2387)* ; 6176GAT(2391)
g2361 and 6177GAT(2389)* 6103GAT(2347)* ; 6181GAT(2392)
g2362 and 6176GAT(2391)* 6175GAT(2390)* ; 6180GAT(2393)
g2363 and 6181GAT(2392)* 6052GAT(2328)* ; 6187GAT(2394)
g2364 and 6181GAT(2392)* 6103GAT(2347)* ; 6185GAT(2395)
g2365 and 6177GAT(2389)* 6181GAT(2392)* ; 6186GAT(2396)
g2366 and 6187GAT(2394)* 6082GAT(2337)* ; 6191GAT(2397)
g2367 and 6186GAT(2396)* 6185GAT(2395)* ; 6190GAT(2398)
g2368 and 6191GAT(2397)* 6026GAT(2315)* ; 6197GAT(2399)
g2369 and 6191GAT(2397)* 6082GAT(2337)* ; 6195GAT(2400)
g2370 and 6187GAT(2394)* 6191GAT(2397)* ; 6196GAT(2401)
g2371 and 6197GAT(2399)* 6058GAT(2325)* ; 6201GAT(2402)
g2372 and 6196GAT(2401)* 6195GAT(2400)* ; 6200GAT(2403)
g2373 and 6201GAT(2402)* 5996GAT(2300)* ; 6207GAT(2404)
g2374 and 6201GAT(2402)* 6058GAT(2325)* ; 6205GAT(2405)
g2375 and 6197GAT(2399)* 6201GAT(2402)* ; 6206GAT(2406)
g2376 and 6207GAT(2404)* 6032GAT(2312)* ; 6211GAT(2407)
g2377 and 6206GAT(2406)* 6205GAT(2405)* ; 6210GAT(2408)
g2378 and 6211GAT(2407)* 5962GAT(2280)* ; 6217GAT(2409)
g2379 and 6211GAT(2407)* 6032GAT(2312)* ; 6215GAT(2410)
g2380 and 6207GAT(2404)* 6211GAT(2407)* ; 6216GAT(2411)
g2381 and 6217GAT(2409)* 6002GAT(2297)* ; 6221GAT(2412)
g2382 and 6216GAT(2411)* 6215GAT(2410)* ; 6220GAT(2413)
g2383 and 6221GAT(2412)* 5919GAT(2261)* ; 6227GAT(2414)
g2384 and 6221GAT(2412)* 6002GAT(2297)* ; 6225GAT(2415)
g2385 and 6217GAT(2409)* 6221GAT(2412)* ; 6226GAT(2416)
g2386 and 6227GAT(2414)* 5968GAT(2277)* ; 6231GAT(2417)
g2387 and 6226GAT(2416)* 6225GAT(2415)* ; 6230GAT(2418)
g2388 and 6231GAT(2417)* 5873GAT(2241)* ; 6237GAT(2419)
g2389 and 6231GAT(2417)* 5968GAT(2277)* ; 6235GAT(2420)
g2390 and 6227GAT(2414)* 6231GAT(2417)* ; 6236GAT(2421)
g2391 and 6237GAT(2419)* 5925GAT(2258)* ; 6241GAT(2422)
g2392 and 6236GAT(2421)* 6235GAT(2420)* ; 6240GAT(2423)
g2393 and 6241GAT(2422)* 5825GAT(2218)* ; 6247GAT(2424)
g2394 and 6241GAT(2422)* 5925GAT(2258)* ; 6245GAT(2425)
g2395 and 6237GAT(2419)* 6241GAT(2422)* ; 6246GAT(2426)
g2396 and 6247GAT(2424)* 5879GAT(2238)* ; 6251GAT(2427)
g2397 and 6246GAT(2426)* 6245GAT(2425)* ; 6250GAT(2428)
g2398 and 6251GAT(2427)* 5776GAT(2195)* ; 6257GAT(2429)
g2399 and 6251GAT(2427)* 5879GAT(2238)* ; 6255GAT(2430)
g2400 and 6247GAT(2424)* 6251GAT(2427)* ; 6256GAT(2431)
g2401 and 6257GAT(2429)* 5831GAT(2215)* ; 6261GAT(2432)
g2402 and 6256GAT(2431)* 6255GAT(2430)* ; 6260GAT(2433)
g2403 and 6261GAT(2432)* 5721GAT(2170)* ; 6267GAT(2434)
g2404 and 6261GAT(2432)* 5831GAT(2215)* ; 6265GAT(2435)
g2405 and 6257GAT(2429)* 6261GAT(2432)* ; 6266GAT(2436)
g2406 and 6267GAT(2434)* 5782GAT(2192)* ; 6271GAT(2437)
g2407 and 6266GAT(2436)* 6265GAT(2435)* ; 6270GAT(2438)
g2408 and 6271GAT(2437)* 5666GAT(2138)* ; 6277GAT(2439)
g2409 and 6271GAT(2437)* 5782GAT(2192)* ; 6275GAT(2440)
g2410 and 6267GAT(2434)* 6271GAT(2437)* ; 6276GAT(2441)
g2411 and 6277GAT(2439)* 5727GAT(2167)* ; 6281GAT(2442)
g2412 and 6276GAT(2441)* 6275GAT(2440)* ; 6280GAT(2443)
g2413 and 6281GAT(2442)* 5602GAT(2110)* ; 6287GAT(2444)
g2414 and 6281GAT(2442)* 5727GAT(2167)* ; 6285GAT(2445)
g2415 and 6277GAT(2439)* 6281GAT(2442)* ; 6286GAT(2446)
g2416 and 6286GAT(2446)* 6285GAT(2445)* ; 6288GAT(2447)
g2417 not 1263GAT(47) ; 1263GAT(47)*
g2418 not 1367GAT(288) ; 1367GAT(288)*
g2419 not 1215GAT(63) ; 1215GAT(63)*
g2420 not 1363GAT(289) ; 1363GAT(289)*
g2421 not 1167GAT(79) ; 1167GAT(79)*
g2422 not 1359GAT(290) ; 1359GAT(290)*
g2423 not 1119GAT(95) ; 1119GAT(95)*
g2424 not 1355GAT(291) ; 1355GAT(291)*
g2425 not 1071GAT(111) ; 1071GAT(111)*
g2426 not 1351GAT(292) ; 1351GAT(292)*
g2427 not 1023GAT(127) ; 1023GAT(127)*
g2428 not 1347GAT(293) ; 1347GAT(293)*
g2429 not 975GAT(143) ; 975GAT(143)*
g2430 not 1343GAT(294) ; 1343GAT(294)*
g2431 not 927GAT(159) ; 927GAT(159)*
g2432 not 1339GAT(295) ; 1339GAT(295)*
g2433 not 879GAT(175) ; 879GAT(175)*
g2434 not 1335GAT(296) ; 1335GAT(296)*
g2435 not 831GAT(191) ; 831GAT(191)*
g2436 not 1331GAT(297) ; 1331GAT(297)*
g2437 not 783GAT(207) ; 783GAT(207)*
g2438 not 1327GAT(298) ; 1327GAT(298)*
g2439 not 735GAT(223) ; 735GAT(223)*
g2440 not 1323GAT(299) ; 1323GAT(299)*
g2441 not 687GAT(239) ; 687GAT(239)*
g2442 not 1319GAT(300) ; 1319GAT(300)*
g2443 not 639GAT(255) ; 639GAT(255)*
g2444 not 1315GAT(301) ; 1315GAT(301)*
g2445 not 591GAT(271) ; 591GAT(271)*
g2446 not 1311GAT(302) ; 1311GAT(302)*
g2447 not 1399GAT(304) ; 1399GAT(304)*
g2448 not 1400GAT(303) ; 1400GAT(303)*
g2449 not 1397GAT(306) ; 1397GAT(306)*
g2450 not 1398GAT(305) ; 1398GAT(305)*
g2451 not 1395GAT(308) ; 1395GAT(308)*
g2452 not 1396GAT(307) ; 1396GAT(307)*
g2453 not 1393GAT(310) ; 1393GAT(310)*
g2454 not 1394GAT(309) ; 1394GAT(309)*
g2455 not 1391GAT(312) ; 1391GAT(312)*
g2456 not 1392GAT(311) ; 1392GAT(311)*
g2457 not 1389GAT(314) ; 1389GAT(314)*
g2458 not 1390GAT(313) ; 1390GAT(313)*
g2459 not 1387GAT(316) ; 1387GAT(316)*
g2460 not 1388GAT(315) ; 1388GAT(315)*
g2461 not 1385GAT(318) ; 1385GAT(318)*
g2462 not 1386GAT(317) ; 1386GAT(317)*
g2463 not 1383GAT(320) ; 1383GAT(320)*
g2464 not 1384GAT(319) ; 1384GAT(319)*
g2465 not 1381GAT(322) ; 1381GAT(322)*
g2466 not 1382GAT(321) ; 1382GAT(321)*
g2467 not 1379GAT(324) ; 1379GAT(324)*
g2468 not 1380GAT(323) ; 1380GAT(323)*
g2469 not 1377GAT(326) ; 1377GAT(326)*
g2470 not 1378GAT(325) ; 1378GAT(325)*
g2471 not 1375GAT(328) ; 1375GAT(328)*
g2472 not 1376GAT(327) ; 1376GAT(327)*
g2473 not 1373GAT(330) ; 1373GAT(330)*
g2474 not 1374GAT(329) ; 1374GAT(329)*
g2475 not 1371GAT(332) ; 1371GAT(332)*
g2476 not 1372GAT(331) ; 1372GAT(331)*
g2477 not 1443GAT(333) ; 1443GAT(333)*
g2478 not 1218GAT(62) ; 1218GAT(62)*
g2479 not 1440GAT(334) ; 1440GAT(334)*
g2480 not 1170GAT(78) ; 1170GAT(78)*
g2481 not 1437GAT(335) ; 1437GAT(335)*
g2482 not 1122GAT(94) ; 1122GAT(94)*
g2483 not 1434GAT(336) ; 1434GAT(336)*
g2484 not 1074GAT(110) ; 1074GAT(110)*
g2485 not 1431GAT(337) ; 1431GAT(337)*
g2486 not 1026GAT(126) ; 1026GAT(126)*
g2487 not 1428GAT(338) ; 1428GAT(338)*
g2488 not 978GAT(142) ; 978GAT(142)*
g2489 not 1425GAT(339) ; 1425GAT(339)*
g2490 not 930GAT(158) ; 930GAT(158)*
g2491 not 1422GAT(340) ; 1422GAT(340)*
g2492 not 882GAT(174) ; 882GAT(174)*
g2493 not 1419GAT(341) ; 1419GAT(341)*
g2494 not 834GAT(190) ; 834GAT(190)*
g2495 not 1416GAT(342) ; 1416GAT(342)*
g2496 not 786GAT(206) ; 786GAT(206)*
g2497 not 1413GAT(343) ; 1413GAT(343)*
g2498 not 738GAT(222) ; 738GAT(222)*
g2499 not 1410GAT(344) ; 1410GAT(344)*
g2500 not 690GAT(238) ; 690GAT(238)*
g2501 not 1407GAT(345) ; 1407GAT(345)*
g2502 not 642GAT(254) ; 642GAT(254)*
g2503 not 1404GAT(346) ; 1404GAT(346)*
g2504 not 594GAT(270) ; 594GAT(270)*
g2505 not 1401GAT(347) ; 1401GAT(347)*
g2506 not 546GAT(286) ; 546GAT(286)*
g2507 not 1502GAT(348) ; 1502GAT(348)*
g2508 not 1498GAT(349) ; 1498GAT(349)*
g2509 not 1494GAT(350) ; 1494GAT(350)*
g2510 not 1490GAT(351) ; 1490GAT(351)*
g2511 not 1486GAT(352) ; 1486GAT(352)*
g2512 not 1482GAT(353) ; 1482GAT(353)*
g2513 not 1478GAT(354) ; 1478GAT(354)*
g2514 not 1474GAT(355) ; 1474GAT(355)*
g2515 not 1470GAT(356) ; 1470GAT(356)*
g2516 not 1466GAT(357) ; 1466GAT(357)*
g2517 not 1462GAT(358) ; 1462GAT(358)*
g2518 not 1458GAT(359) ; 1458GAT(359)*
g2519 not 1454GAT(360) ; 1454GAT(360)*
g2520 not 1450GAT(361) ; 1450GAT(361)*
g2521 not 1446GAT(362) ; 1446GAT(362)*
g2522 not 1266GAT(46) ; 1266GAT(46)*
g2523 not 1578GAT(363) ; 1578GAT(363)*
g2524 not 1576GAT(364) ; 1576GAT(364)*
g2525 not 1577GAT(365) ; 1577GAT(365)*
g2526 not 1571GAT(367) ; 1571GAT(367)*
g2527 not 1572GAT(368) ; 1572GAT(368)*
g2528 not 1566GAT(370) ; 1566GAT(370)*
g2529 not 1567GAT(371) ; 1567GAT(371)*
g2530 not 1561GAT(373) ; 1561GAT(373)*
g2531 not 1562GAT(374) ; 1562GAT(374)*
g2532 not 1556GAT(376) ; 1556GAT(376)*
g2533 not 1557GAT(377) ; 1557GAT(377)*
g2534 not 1551GAT(379) ; 1551GAT(379)*
g2535 not 1552GAT(380) ; 1552GAT(380)*
g2536 not 1546GAT(382) ; 1546GAT(382)*
g2537 not 1547GAT(383) ; 1547GAT(383)*
g2538 not 1541GAT(385) ; 1541GAT(385)*
g2539 not 1542GAT(386) ; 1542GAT(386)*
g2540 not 1536GAT(388) ; 1536GAT(388)*
g2541 not 1537GAT(389) ; 1537GAT(389)*
g2542 not 1531GAT(391) ; 1531GAT(391)*
g2543 not 1532GAT(392) ; 1532GAT(392)*
g2544 not 1526GAT(394) ; 1526GAT(394)*
g2545 not 1527GAT(395) ; 1527GAT(395)*
g2546 not 1521GAT(397) ; 1521GAT(397)*
g2547 not 1522GAT(398) ; 1522GAT(398)*
g2548 not 1516GAT(400) ; 1516GAT(400)*
g2549 not 1517GAT(401) ; 1517GAT(401)*
g2550 not 1511GAT(403) ; 1511GAT(403)*
g2551 not 1512GAT(404) ; 1512GAT(404)*
g2552 not 1506GAT(406) ; 1506GAT(406)*
g2553 not 1507GAT(407) ; 1507GAT(407)*
g2554 not 1624GAT(408) ; 1624GAT(408)*
g2555 not 1621GAT(409) ; 1621GAT(409)*
g2556 not 1573GAT(366) ; 1573GAT(366)*
g2557 not 1618GAT(410) ; 1618GAT(410)*
g2558 not 1568GAT(369) ; 1568GAT(369)*
g2559 not 1615GAT(411) ; 1615GAT(411)*
g2560 not 1563GAT(372) ; 1563GAT(372)*
g2561 not 1612GAT(412) ; 1612GAT(412)*
g2562 not 1558GAT(375) ; 1558GAT(375)*
g2563 not 1609GAT(413) ; 1609GAT(413)*
g2564 not 1553GAT(378) ; 1553GAT(378)*
g2565 not 1606GAT(414) ; 1606GAT(414)*
g2566 not 1548GAT(381) ; 1548GAT(381)*
g2567 not 1603GAT(415) ; 1603GAT(415)*
g2568 not 1543GAT(384) ; 1543GAT(384)*
g2569 not 1600GAT(416) ; 1600GAT(416)*
g2570 not 1538GAT(387) ; 1538GAT(387)*
g2571 not 1597GAT(417) ; 1597GAT(417)*
g2572 not 1533GAT(390) ; 1533GAT(390)*
g2573 not 1594GAT(418) ; 1594GAT(418)*
g2574 not 1528GAT(393) ; 1528GAT(393)*
g2575 not 1591GAT(419) ; 1591GAT(419)*
g2576 not 1523GAT(396) ; 1523GAT(396)*
g2577 not 1588GAT(420) ; 1588GAT(420)*
g2578 not 1518GAT(399) ; 1518GAT(399)*
g2579 not 1585GAT(421) ; 1585GAT(421)*
g2580 not 1513GAT(402) ; 1513GAT(402)*
g2581 not 1582GAT(422) ; 1582GAT(422)*
g2582 not 1508GAT(405) ; 1508GAT(405)*
g2583 not 1684GAT(424) ; 1684GAT(424)*
g2584 not 1685GAT(425) ; 1685GAT(425)*
g2585 not 1680GAT(426) ; 1680GAT(426)*
g2586 not 1676GAT(427) ; 1676GAT(427)*
g2587 not 1672GAT(428) ; 1672GAT(428)*
g2588 not 1668GAT(429) ; 1668GAT(429)*
g2589 not 1664GAT(430) ; 1664GAT(430)*
g2590 not 1660GAT(431) ; 1660GAT(431)*
g2591 not 1656GAT(432) ; 1656GAT(432)*
g2592 not 1652GAT(433) ; 1652GAT(433)*
g2593 not 1648GAT(434) ; 1648GAT(434)*
g2594 not 1644GAT(435) ; 1644GAT(435)*
g2595 not 1640GAT(436) ; 1640GAT(436)*
g2596 not 1636GAT(437) ; 1636GAT(437)*
g2597 not 1632GAT(438) ; 1632GAT(438)*
g2598 not 1628GAT(439) ; 1628GAT(439)*
g2599 not 1712GAT(441) ; 1712GAT(441)*
g2600 not 1713GAT(442) ; 1713GAT(442)*
g2601 not 1714GAT(440) ; 1714GAT(440)*
g2602 not 1221GAT(61) ; 1221GAT(61)*
g2603 not 1710GAT(443) ; 1710GAT(443)*
g2604 not 1711GAT(444) ; 1711GAT(444)*
g2605 not 1708GAT(445) ; 1708GAT(445)*
g2606 not 1709GAT(446) ; 1709GAT(446)*
g2607 not 1706GAT(447) ; 1706GAT(447)*
g2608 not 1707GAT(448) ; 1707GAT(448)*
g2609 not 1704GAT(449) ; 1704GAT(449)*
g2610 not 1705GAT(450) ; 1705GAT(450)*
g2611 not 1702GAT(451) ; 1702GAT(451)*
g2612 not 1703GAT(452) ; 1703GAT(452)*
g2613 not 1700GAT(453) ; 1700GAT(453)*
g2614 not 1701GAT(454) ; 1701GAT(454)*
g2615 not 1698GAT(455) ; 1698GAT(455)*
g2616 not 1699GAT(456) ; 1699GAT(456)*
g2617 not 1696GAT(457) ; 1696GAT(457)*
g2618 not 1697GAT(458) ; 1697GAT(458)*
g2619 not 1694GAT(459) ; 1694GAT(459)*
g2620 not 1695GAT(460) ; 1695GAT(460)*
g2621 not 1692GAT(461) ; 1692GAT(461)*
g2622 not 1693GAT(462) ; 1693GAT(462)*
g2623 not 1690GAT(463) ; 1690GAT(463)*
g2624 not 1691GAT(464) ; 1691GAT(464)*
g2625 not 1688GAT(465) ; 1688GAT(465)*
g2626 not 1689GAT(466) ; 1689GAT(466)*
g2627 not 1686GAT(467) ; 1686GAT(467)*
g2628 not 1687GAT(468) ; 1687GAT(468)*
g2629 not 1759GAT(470) ; 1759GAT(470)*
g2630 not 1756GAT(469) ; 1756GAT(469)*
g2631 not 1173GAT(77) ; 1173GAT(77)*
g2632 not 1753GAT(471) ; 1753GAT(471)*
g2633 not 1125GAT(93) ; 1125GAT(93)*
g2634 not 1750GAT(472) ; 1750GAT(472)*
g2635 not 1077GAT(109) ; 1077GAT(109)*
g2636 not 1747GAT(473) ; 1747GAT(473)*
g2637 not 1029GAT(125) ; 1029GAT(125)*
g2638 not 1744GAT(474) ; 1744GAT(474)*
g2639 not 981GAT(141) ; 981GAT(141)*
g2640 not 1741GAT(475) ; 1741GAT(475)*
g2641 not 933GAT(157) ; 933GAT(157)*
g2642 not 1738GAT(476) ; 1738GAT(476)*
g2643 not 885GAT(173) ; 885GAT(173)*
g2644 not 1735GAT(477) ; 1735GAT(477)*
g2645 not 837GAT(189) ; 837GAT(189)*
g2646 not 1732GAT(478) ; 1732GAT(478)*
g2647 not 789GAT(205) ; 789GAT(205)*
g2648 not 1729GAT(479) ; 1729GAT(479)*
g2649 not 741GAT(221) ; 741GAT(221)*
g2650 not 1726GAT(480) ; 1726GAT(480)*
g2651 not 693GAT(237) ; 693GAT(237)*
g2652 not 1723GAT(481) ; 1723GAT(481)*
g2653 not 645GAT(253) ; 645GAT(253)*
g2654 not 1720GAT(482) ; 1720GAT(482)*
g2655 not 597GAT(269) ; 597GAT(269)*
g2656 not 1717GAT(483) ; 1717GAT(483)*
g2657 not 549GAT(285) ; 549GAT(285)*
g2658 not 1269GAT(45) ; 1269GAT(45)*
g2659 not 1821GAT(484) ; 1821GAT(484)*
g2660 not 1819GAT(485) ; 1819GAT(485)*
g2661 not 1820GAT(486) ; 1820GAT(486)*
g2662 not 1815GAT(487) ; 1815GAT(487)*
g2663 not 1811GAT(488) ; 1811GAT(488)*
g2664 not 1807GAT(489) ; 1807GAT(489)*
g2665 not 1803GAT(490) ; 1803GAT(490)*
g2666 not 1799GAT(491) ; 1799GAT(491)*
g2667 not 1795GAT(492) ; 1795GAT(492)*
g2668 not 1791GAT(493) ; 1791GAT(493)*
g2669 not 1787GAT(494) ; 1787GAT(494)*
g2670 not 1783GAT(495) ; 1783GAT(495)*
g2671 not 1779GAT(496) ; 1779GAT(496)*
g2672 not 1775GAT(497) ; 1775GAT(497)*
g2673 not 1771GAT(498) ; 1771GAT(498)*
g2674 not 1767GAT(499) ; 1767GAT(499)*
g2675 not 1763GAT(500) ; 1763GAT(500)*
g2676 not 1897GAT(501) ; 1897GAT(501)*
g2677 not 1894GAT(502) ; 1894GAT(502)*
g2678 not 1891GAT(504) ; 1891GAT(504)*
g2679 not 1889GAT(503) ; 1889GAT(503)*
g2680 not 1890GAT(506) ; 1890GAT(506)*
g2681 not 1884GAT(505) ; 1884GAT(505)*
g2682 not 1885GAT(509) ; 1885GAT(509)*
g2683 not 1879GAT(508) ; 1879GAT(508)*
g2684 not 1880GAT(512) ; 1880GAT(512)*
g2685 not 1874GAT(511) ; 1874GAT(511)*
g2686 not 1875GAT(515) ; 1875GAT(515)*
g2687 not 1869GAT(514) ; 1869GAT(514)*
g2688 not 1870GAT(518) ; 1870GAT(518)*
g2689 not 1864GAT(517) ; 1864GAT(517)*
g2690 not 1865GAT(521) ; 1865GAT(521)*
g2691 not 1859GAT(520) ; 1859GAT(520)*
g2692 not 1860GAT(524) ; 1860GAT(524)*
g2693 not 1854GAT(523) ; 1854GAT(523)*
g2694 not 1855GAT(527) ; 1855GAT(527)*
g2695 not 1849GAT(526) ; 1849GAT(526)*
g2696 not 1850GAT(530) ; 1850GAT(530)*
g2697 not 1844GAT(529) ; 1844GAT(529)*
g2698 not 1845GAT(533) ; 1845GAT(533)*
g2699 not 1839GAT(532) ; 1839GAT(532)*
g2700 not 1840GAT(536) ; 1840GAT(536)*
g2701 not 1834GAT(535) ; 1834GAT(535)*
g2702 not 1835GAT(539) ; 1835GAT(539)*
g2703 not 1829GAT(538) ; 1829GAT(538)*
g2704 not 1830GAT(542) ; 1830GAT(542)*
g2705 not 1824GAT(541) ; 1824GAT(541)*
g2706 not 1825GAT(544) ; 1825GAT(544)*
g2707 not 1945GAT(545) ; 1945GAT(545)*
g2708 not 1946GAT(546) ; 1946GAT(546)*
g2709 not 1941GAT(547) ; 1941GAT(547)*
g2710 not 1938GAT(548) ; 1938GAT(548)*
g2711 not 1886GAT(507) ; 1886GAT(507)*
g2712 not 1935GAT(549) ; 1935GAT(549)*
g2713 not 1881GAT(510) ; 1881GAT(510)*
g2714 not 1932GAT(550) ; 1932GAT(550)*
g2715 not 1876GAT(513) ; 1876GAT(513)*
g2716 not 1929GAT(551) ; 1929GAT(551)*
g2717 not 1871GAT(516) ; 1871GAT(516)*
g2718 not 1926GAT(552) ; 1926GAT(552)*
g2719 not 1866GAT(519) ; 1866GAT(519)*
g2720 not 1923GAT(553) ; 1923GAT(553)*
g2721 not 1861GAT(522) ; 1861GAT(522)*
g2722 not 1920GAT(554) ; 1920GAT(554)*
g2723 not 1856GAT(525) ; 1856GAT(525)*
g2724 not 1917GAT(555) ; 1917GAT(555)*
g2725 not 1851GAT(528) ; 1851GAT(528)*
g2726 not 1914GAT(556) ; 1914GAT(556)*
g2727 not 1846GAT(531) ; 1846GAT(531)*
g2728 not 1911GAT(557) ; 1911GAT(557)*
g2729 not 1841GAT(534) ; 1841GAT(534)*
g2730 not 1908GAT(558) ; 1908GAT(558)*
g2731 not 1836GAT(537) ; 1836GAT(537)*
g2732 not 1905GAT(559) ; 1905GAT(559)*
g2733 not 1831GAT(540) ; 1831GAT(540)*
g2734 not 1902GAT(560) ; 1902GAT(560)*
g2735 not 1826GAT(543) ; 1826GAT(543)*
g2736 not 1999GAT(563) ; 1999GAT(563)*
g2737 not 2000GAT(564) ; 2000GAT(564)*
g2738 not 1995GAT(565) ; 1995GAT(565)*
g2739 not 2001GAT(562) ; 2001GAT(562)*
g2740 not 1224GAT(60) ; 1224GAT(60)*
g2741 not 1991GAT(566) ; 1991GAT(566)*
g2742 not 1987GAT(567) ; 1987GAT(567)*
g2743 not 1983GAT(568) ; 1983GAT(568)*
g2744 not 1979GAT(569) ; 1979GAT(569)*
g2745 not 1975GAT(570) ; 1975GAT(570)*
g2746 not 1971GAT(571) ; 1971GAT(571)*
g2747 not 1967GAT(572) ; 1967GAT(572)*
g2748 not 1963GAT(573) ; 1963GAT(573)*
g2749 not 1959GAT(574) ; 1959GAT(574)*
g2750 not 1955GAT(575) ; 1955GAT(575)*
g2751 not 1951GAT(576) ; 1951GAT(576)*
g2752 not 1947GAT(577) ; 1947GAT(577)*
g2753 not 2033GAT(580) ; 2033GAT(580)*
g2754 not 2028GAT(579) ; 2028GAT(579)*
g2755 not 2029GAT(582) ; 2029GAT(582)*
g2756 not 2026GAT(581) ; 2026GAT(581)*
g2757 not 2027GAT(584) ; 2027GAT(584)*
g2758 not 2030GAT(578) ; 2030GAT(578)*
g2759 not 1176GAT(76) ; 1176GAT(76)*
g2760 not 2024GAT(583) ; 2024GAT(583)*
g2761 not 2025GAT(586) ; 2025GAT(586)*
g2762 not 2022GAT(585) ; 2022GAT(585)*
g2763 not 2023GAT(588) ; 2023GAT(588)*
g2764 not 2020GAT(587) ; 2020GAT(587)*
g2765 not 2021GAT(590) ; 2021GAT(590)*
g2766 not 2018GAT(589) ; 2018GAT(589)*
g2767 not 2019GAT(592) ; 2019GAT(592)*
g2768 not 2016GAT(591) ; 2016GAT(591)*
g2769 not 2017GAT(594) ; 2017GAT(594)*
g2770 not 2014GAT(593) ; 2014GAT(593)*
g2771 not 2015GAT(596) ; 2015GAT(596)*
g2772 not 2012GAT(595) ; 2012GAT(595)*
g2773 not 2013GAT(598) ; 2013GAT(598)*
g2774 not 2010GAT(597) ; 2010GAT(597)*
g2775 not 2011GAT(600) ; 2011GAT(600)*
g2776 not 2008GAT(599) ; 2008GAT(599)*
g2777 not 2009GAT(602) ; 2009GAT(602)*
g2778 not 2006GAT(601) ; 2006GAT(601)*
g2779 not 2007GAT(604) ; 2007GAT(604)*
g2780 not 2004GAT(603) ; 2004GAT(603)*
g2781 not 2005GAT(605) ; 2005GAT(605)*
g2782 not 1272GAT(44) ; 1272GAT(44)*
g2783 not 2082GAT(606) ; 2082GAT(606)*
g2784 not 2080GAT(607) ; 2080GAT(607)*
g2785 not 2081GAT(609) ; 2081GAT(609)*
g2786 not 2076GAT(611) ; 2076GAT(611)*
g2787 not 2073GAT(608) ; 2073GAT(608)*
g2788 not 1128GAT(92) ; 1128GAT(92)*
g2789 not 2070GAT(610) ; 2070GAT(610)*
g2790 not 1080GAT(108) ; 1080GAT(108)*
g2791 not 2067GAT(612) ; 2067GAT(612)*
g2792 not 1032GAT(124) ; 1032GAT(124)*
g2793 not 2064GAT(613) ; 2064GAT(613)*
g2794 not 984GAT(140) ; 984GAT(140)*
g2795 not 2061GAT(614) ; 2061GAT(614)*
g2796 not 936GAT(156) ; 936GAT(156)*
g2797 not 2058GAT(615) ; 2058GAT(615)*
g2798 not 888GAT(172) ; 888GAT(172)*
g2799 not 2055GAT(616) ; 2055GAT(616)*
g2800 not 840GAT(188) ; 840GAT(188)*
g2801 not 2052GAT(617) ; 2052GAT(617)*
g2802 not 792GAT(204) ; 792GAT(204)*
g2803 not 2049GAT(618) ; 2049GAT(618)*
g2804 not 744GAT(220) ; 744GAT(220)*
g2805 not 2046GAT(619) ; 2046GAT(619)*
g2806 not 696GAT(236) ; 696GAT(236)*
g2807 not 2043GAT(620) ; 2043GAT(620)*
g2808 not 648GAT(252) ; 648GAT(252)*
g2809 not 2040GAT(621) ; 2040GAT(621)*
g2810 not 600GAT(268) ; 600GAT(268)*
g2811 not 2037GAT(622) ; 2037GAT(622)*
g2812 not 552GAT(284) ; 552GAT(284)*
g2813 not 2145GAT(623) ; 2145GAT(623)*
g2814 not 2142GAT(624) ; 2142GAT(624)*
g2815 not 2139GAT(625) ; 2139GAT(625)*
g2816 not 2137GAT(626) ; 2137GAT(626)*
g2817 not 2138GAT(627) ; 2138GAT(627)*
g2818 not 2133GAT(628) ; 2133GAT(628)*
g2819 not 2129GAT(629) ; 2129GAT(629)*
g2820 not 2125GAT(630) ; 2125GAT(630)*
g2821 not 2121GAT(631) ; 2121GAT(631)*
g2822 not 2117GAT(632) ; 2117GAT(632)*
g2823 not 2113GAT(633) ; 2113GAT(633)*
g2824 not 2109GAT(634) ; 2109GAT(634)*
g2825 not 2105GAT(635) ; 2105GAT(635)*
g2826 not 2101GAT(636) ; 2101GAT(636)*
g2827 not 2097GAT(637) ; 2097GAT(637)*
g2828 not 2093GAT(638) ; 2093GAT(638)*
g2829 not 2089GAT(639) ; 2089GAT(639)*
g2830 not 2085GAT(640) ; 2085GAT(640)*
g2831 not 2221GAT(641) ; 2221GAT(641)*
g2832 not 2222GAT(642) ; 2222GAT(642)*
g2833 not 2217GAT(643) ; 2217GAT(643)*
g2834 not 2214GAT(644) ; 2214GAT(644)*
g2835 not 2211GAT(647) ; 2211GAT(647)*
g2836 not 2209GAT(645) ; 2209GAT(645)*
g2837 not 2210GAT(649) ; 2210GAT(649)*
g2838 not 2204GAT(646) ; 2204GAT(646)*
g2839 not 2205GAT(652) ; 2205GAT(652)*
g2840 not 2199GAT(648) ; 2199GAT(648)*
g2841 not 2200GAT(655) ; 2200GAT(655)*
g2842 not 2194GAT(651) ; 2194GAT(651)*
g2843 not 2195GAT(658) ; 2195GAT(658)*
g2844 not 2189GAT(654) ; 2189GAT(654)*
g2845 not 2190GAT(661) ; 2190GAT(661)*
g2846 not 2184GAT(657) ; 2184GAT(657)*
g2847 not 2185GAT(664) ; 2185GAT(664)*
g2848 not 2179GAT(660) ; 2179GAT(660)*
g2849 not 2180GAT(667) ; 2180GAT(667)*
g2850 not 2174GAT(663) ; 2174GAT(663)*
g2851 not 2175GAT(670) ; 2175GAT(670)*
g2852 not 2169GAT(666) ; 2169GAT(666)*
g2853 not 2170GAT(673) ; 2170GAT(673)*
g2854 not 2164GAT(669) ; 2164GAT(669)*
g2855 not 2165GAT(676) ; 2165GAT(676)*
g2856 not 2159GAT(672) ; 2159GAT(672)*
g2857 not 2160GAT(679) ; 2160GAT(679)*
g2858 not 2154GAT(675) ; 2154GAT(675)*
g2859 not 2155GAT(681) ; 2155GAT(681)*
g2860 not 2149GAT(678) ; 2149GAT(678)*
g2861 not 2150GAT(683) ; 2150GAT(683)*
g2862 not 2264GAT(685) ; 2264GAT(685)*
g2863 not 2265GAT(686) ; 2265GAT(686)*
g2864 not 2260GAT(687) ; 2260GAT(687)*
g2865 not 2266GAT(684) ; 2266GAT(684)*
g2866 not 1227GAT(59) ; 1227GAT(59)*
g2867 not 2257GAT(688) ; 2257GAT(688)*
g2868 not 2206GAT(650) ; 2206GAT(650)*
g2869 not 2254GAT(689) ; 2254GAT(689)*
g2870 not 2201GAT(653) ; 2201GAT(653)*
g2871 not 2251GAT(690) ; 2251GAT(690)*
g2872 not 2196GAT(656) ; 2196GAT(656)*
g2873 not 2248GAT(691) ; 2248GAT(691)*
g2874 not 2191GAT(659) ; 2191GAT(659)*
g2875 not 2245GAT(692) ; 2245GAT(692)*
g2876 not 2186GAT(662) ; 2186GAT(662)*
g2877 not 2242GAT(693) ; 2242GAT(693)*
g2878 not 2181GAT(665) ; 2181GAT(665)*
g2879 not 2239GAT(694) ; 2239GAT(694)*
g2880 not 2176GAT(668) ; 2176GAT(668)*
g2881 not 2236GAT(695) ; 2236GAT(695)*
g2882 not 2171GAT(671) ; 2171GAT(671)*
g2883 not 2233GAT(696) ; 2233GAT(696)*
g2884 not 2166GAT(674) ; 2166GAT(674)*
g2885 not 2230GAT(697) ; 2230GAT(697)*
g2886 not 2161GAT(677) ; 2161GAT(677)*
g2887 not 2227GAT(698) ; 2227GAT(698)*
g2888 not 2156GAT(680) ; 2156GAT(680)*
g2889 not 2224GAT(699) ; 2224GAT(699)*
g2890 not 2151GAT(682) ; 2151GAT(682)*
g2891 not 2322GAT(703) ; 2322GAT(703)*
g2892 not 2317GAT(702) ; 2317GAT(702)*
g2893 not 2318GAT(704) ; 2318GAT(704)*
g2894 not 2313GAT(705) ; 2313GAT(705)*
g2895 not 2309GAT(706) ; 2309GAT(706)*
g2896 not 2319GAT(701) ; 2319GAT(701)*
g2897 not 1179GAT(75) ; 1179GAT(75)*
g2898 not 2305GAT(707) ; 2305GAT(707)*
g2899 not 2301GAT(708) ; 2301GAT(708)*
g2900 not 2297GAT(709) ; 2297GAT(709)*
g2901 not 2293GAT(710) ; 2293GAT(710)*
g2902 not 2289GAT(711) ; 2289GAT(711)*
g2903 not 2285GAT(712) ; 2285GAT(712)*
g2904 not 2281GAT(713) ; 2281GAT(713)*
g2905 not 2277GAT(714) ; 2277GAT(714)*
g2906 not 2273GAT(715) ; 2273GAT(715)*
g2907 not 2269GAT(716) ; 2269GAT(716)*
g2908 not 1275GAT(43) ; 1275GAT(43)*
g2909 not 2359GAT(717) ; 2359GAT(717)*
g2910 not 2357GAT(718) ; 2357GAT(718)*
g2911 not 2358GAT(721) ; 2358GAT(721)*
g2912 not 2353GAT(723) ; 2353GAT(723)*
g2913 not 2348GAT(720) ; 2348GAT(720)*
g2914 not 2349GAT(725) ; 2349GAT(725)*
g2915 not 2346GAT(722) ; 2346GAT(722)*
g2916 not 2347GAT(727) ; 2347GAT(727)*
g2917 not 2344GAT(724) ; 2344GAT(724)*
g2918 not 2345GAT(729) ; 2345GAT(729)*
g2919 not 2350GAT(719) ; 2350GAT(719)*
g2920 not 1131GAT(91) ; 1131GAT(91)*
g2921 not 2342GAT(726) ; 2342GAT(726)*
g2922 not 2343GAT(731) ; 2343GAT(731)*
g2923 not 2340GAT(728) ; 2340GAT(728)*
g2924 not 2341GAT(733) ; 2341GAT(733)*
g2925 not 2338GAT(730) ; 2338GAT(730)*
g2926 not 2339GAT(735) ; 2339GAT(735)*
g2927 not 2336GAT(732) ; 2336GAT(732)*
g2928 not 2337GAT(737) ; 2337GAT(737)*
g2929 not 2334GAT(734) ; 2334GAT(734)*
g2930 not 2335GAT(739) ; 2335GAT(739)*
g2931 not 2332GAT(736) ; 2332GAT(736)*
g2932 not 2333GAT(741) ; 2333GAT(741)*
g2933 not 2330GAT(738) ; 2330GAT(738)*
g2934 not 2331GAT(743) ; 2331GAT(743)*
g2935 not 2328GAT(740) ; 2328GAT(740)*
g2936 not 2329GAT(744) ; 2329GAT(744)*
g2937 not 2326GAT(742) ; 2326GAT(742)*
g2938 not 2327GAT(745) ; 2327GAT(745)*
g2939 not 2410GAT(746) ; 2410GAT(746)*
g2940 not 2407GAT(747) ; 2407GAT(747)*
g2941 not 2404GAT(748) ; 2404GAT(748)*
g2942 not 2402GAT(749) ; 2402GAT(749)*
g2943 not 2403GAT(752) ; 2403GAT(752)*
g2944 not 2398GAT(754) ; 2398GAT(754)*
g2945 not 2395GAT(750) ; 2395GAT(750)*
g2946 not 1083GAT(107) ; 1083GAT(107)*
g2947 not 2392GAT(751) ; 2392GAT(751)*
g2948 not 1035GAT(123) ; 1035GAT(123)*
g2949 not 2389GAT(753) ; 2389GAT(753)*
g2950 not 987GAT(139) ; 987GAT(139)*
g2951 not 2386GAT(755) ; 2386GAT(755)*
g2952 not 939GAT(155) ; 939GAT(155)*
g2953 not 2383GAT(756) ; 2383GAT(756)*
g2954 not 891GAT(171) ; 891GAT(171)*
g2955 not 2380GAT(757) ; 2380GAT(757)*
g2956 not 843GAT(187) ; 843GAT(187)*
g2957 not 2377GAT(758) ; 2377GAT(758)*
g2958 not 795GAT(203) ; 795GAT(203)*
g2959 not 2374GAT(759) ; 2374GAT(759)*
g2960 not 747GAT(219) ; 747GAT(219)*
g2961 not 2371GAT(760) ; 2371GAT(760)*
g2962 not 699GAT(235) ; 699GAT(235)*
g2963 not 2368GAT(761) ; 2368GAT(761)*
g2964 not 651GAT(251) ; 651GAT(251)*
g2965 not 2365GAT(762) ; 2365GAT(762)*
g2966 not 603GAT(267) ; 603GAT(267)*
g2967 not 2362GAT(763) ; 2362GAT(763)*
g2968 not 555GAT(283) ; 555GAT(283)*
g2969 not 2474GAT(764) ; 2474GAT(764)*
g2970 not 2475GAT(765) ; 2475GAT(765)*
g2971 not 2470GAT(766) ; 2470GAT(766)*
g2972 not 2467GAT(767) ; 2467GAT(767)*
g2973 not 2464GAT(768) ; 2464GAT(768)*
g2974 not 2462GAT(769) ; 2462GAT(769)*
g2975 not 2463GAT(770) ; 2463GAT(770)*
g2976 not 2458GAT(771) ; 2458GAT(771)*
g2977 not 2454GAT(772) ; 2454GAT(772)*
g2978 not 2450GAT(773) ; 2450GAT(773)*
g2979 not 2446GAT(774) ; 2446GAT(774)*
g2980 not 2442GAT(775) ; 2442GAT(775)*
g2981 not 2438GAT(776) ; 2438GAT(776)*
g2982 not 2434GAT(777) ; 2434GAT(777)*
g2983 not 2430GAT(778) ; 2430GAT(778)*
g2984 not 2426GAT(779) ; 2426GAT(779)*
g2985 not 2422GAT(780) ; 2422GAT(780)*
g2986 not 2418GAT(781) ; 2418GAT(781)*
g2987 not 2414GAT(782) ; 2414GAT(782)*
g2988 not 2543GAT(784) ; 2543GAT(784)*
g2989 not 2544GAT(785) ; 2544GAT(785)*
g2990 not 2539GAT(786) ; 2539GAT(786)*
g2991 not 2536GAT(787) ; 2536GAT(787)*
g2992 not 2533GAT(791) ; 2533GAT(791)*
g2993 not 2531GAT(788) ; 2531GAT(788)*
g2994 not 2532GAT(793) ; 2532GAT(793)*
g2995 not 2545GAT(783) ; 2545GAT(783)*
g2996 not 1230GAT(58) ; 1230GAT(58)*
g2997 not 2526GAT(789) ; 2526GAT(789)*
g2998 not 2527GAT(796) ; 2527GAT(796)*
g2999 not 2521GAT(790) ; 2521GAT(790)*
g3000 not 2522GAT(799) ; 2522GAT(799)*
g3001 not 2516GAT(792) ; 2516GAT(792)*
g3002 not 2517GAT(802) ; 2517GAT(802)*
g3003 not 2511GAT(795) ; 2511GAT(795)*
g3004 not 2512GAT(805) ; 2512GAT(805)*
g3005 not 2506GAT(798) ; 2506GAT(798)*
g3006 not 2507GAT(808) ; 2507GAT(808)*
g3007 not 2501GAT(801) ; 2501GAT(801)*
g3008 not 2502GAT(811) ; 2502GAT(811)*
g3009 not 2496GAT(804) ; 2496GAT(804)*
g3010 not 2497GAT(814) ; 2497GAT(814)*
g3011 not 2491GAT(807) ; 2491GAT(807)*
g3012 not 2492GAT(817) ; 2492GAT(817)*
g3013 not 2486GAT(810) ; 2486GAT(810)*
g3014 not 2487GAT(819) ; 2487GAT(819)*
g3015 not 2481GAT(813) ; 2481GAT(813)*
g3016 not 2482GAT(821) ; 2482GAT(821)*
g3017 not 2476GAT(816) ; 2476GAT(816)*
g3018 not 2477GAT(823) ; 2477GAT(823)*
g3019 not 2591GAT(829) ; 2591GAT(829)*
g3020 not 2586GAT(825) ; 2586GAT(825)*
g3021 not 2587GAT(826) ; 2587GAT(826)*
g3022 not 2582GAT(827) ; 2582GAT(827)*
g3023 not 2588GAT(824) ; 2588GAT(824)*
g3024 not 1182GAT(74) ; 1182GAT(74)*
g3025 not 2579GAT(828) ; 2579GAT(828)*
g3026 not 2528GAT(794) ; 2528GAT(794)*
g3027 not 2576GAT(830) ; 2576GAT(830)*
g3028 not 2523GAT(797) ; 2523GAT(797)*
g3029 not 2573GAT(831) ; 2573GAT(831)*
g3030 not 2518GAT(800) ; 2518GAT(800)*
g3031 not 2570GAT(832) ; 2570GAT(832)*
g3032 not 2513GAT(803) ; 2513GAT(803)*
g3033 not 2567GAT(833) ; 2567GAT(833)*
g3034 not 2508GAT(806) ; 2508GAT(806)*
g3035 not 2564GAT(834) ; 2564GAT(834)*
g3036 not 2503GAT(809) ; 2503GAT(809)*
g3037 not 2561GAT(835) ; 2561GAT(835)*
g3038 not 2498GAT(812) ; 2498GAT(812)*
g3039 not 2558GAT(836) ; 2558GAT(836)*
g3040 not 2493GAT(815) ; 2493GAT(815)*
g3041 not 2555GAT(837) ; 2555GAT(837)*
g3042 not 2488GAT(818) ; 2488GAT(818)*
g3043 not 2552GAT(838) ; 2552GAT(838)*
g3044 not 2483GAT(820) ; 2483GAT(820)*
g3045 not 2549GAT(839) ; 2549GAT(839)*
g3046 not 2478GAT(822) ; 2478GAT(822)*
g3047 not 1278GAT(42) ; 1278GAT(42)*
g3048 not 2650GAT(841) ; 2650GAT(841)*
g3049 not 2648GAT(842) ; 2648GAT(842)*
g3050 not 2649GAT(845) ; 2649GAT(845)*
g3051 not 2644GAT(846) ; 2644GAT(846)*
g3052 not 2639GAT(844) ; 2639GAT(844)*
g3053 not 2640GAT(847) ; 2640GAT(847)*
g3054 not 2635GAT(848) ; 2635GAT(848)*
g3055 not 2631GAT(849) ; 2631GAT(849)*
g3056 not 2627GAT(850) ; 2627GAT(850)*
g3057 not 2641GAT(843) ; 2641GAT(843)*
g3058 not 1134GAT(90) ; 1134GAT(90)*
g3059 not 2623GAT(851) ; 2623GAT(851)*
g3060 not 2619GAT(852) ; 2619GAT(852)*
g3061 not 2615GAT(853) ; 2615GAT(853)*
g3062 not 2611GAT(854) ; 2611GAT(854)*
g3063 not 2607GAT(855) ; 2607GAT(855)*
g3064 not 2603GAT(856) ; 2603GAT(856)*
g3065 not 2599GAT(857) ; 2599GAT(857)*
g3066 not 2595GAT(858) ; 2595GAT(858)*
g3067 not 2690GAT(859) ; 2690GAT(859)*
g3068 not 2687GAT(860) ; 2687GAT(860)*
g3069 not 2684GAT(861) ; 2684GAT(861)*
g3070 not 2682GAT(862) ; 2682GAT(862)*
g3071 not 2683GAT(866) ; 2683GAT(866)*
g3072 not 2678GAT(868) ; 2678GAT(868)*
g3073 not 2673GAT(864) ; 2673GAT(864)*
g3074 not 2674GAT(870) ; 2674GAT(870)*
g3075 not 2671GAT(865) ; 2671GAT(865)*
g3076 not 2672GAT(872) ; 2672GAT(872)*
g3077 not 2669GAT(867) ; 2669GAT(867)*
g3078 not 2670GAT(874) ; 2670GAT(874)*
g3079 not 2667GAT(869) ; 2667GAT(869)*
g3080 not 2668GAT(876) ; 2668GAT(876)*
g3081 not 2675GAT(863) ; 2675GAT(863)*
g3082 not 1086GAT(106) ; 1086GAT(106)*
g3083 not 2665GAT(871) ; 2665GAT(871)*
g3084 not 2666GAT(878) ; 2666GAT(878)*
g3085 not 2663GAT(873) ; 2663GAT(873)*
g3086 not 2664GAT(880) ; 2664GAT(880)*
g3087 not 2661GAT(875) ; 2661GAT(875)*
g3088 not 2662GAT(882) ; 2662GAT(882)*
g3089 not 2659GAT(877) ; 2659GAT(877)*
g3090 not 2660GAT(884) ; 2660GAT(884)*
g3091 not 2657GAT(879) ; 2657GAT(879)*
g3092 not 2658GAT(885) ; 2658GAT(885)*
g3093 not 2655GAT(881) ; 2655GAT(881)*
g3094 not 2656GAT(886) ; 2656GAT(886)*
g3095 not 2653GAT(883) ; 2653GAT(883)*
g3096 not 2654GAT(887) ; 2654GAT(887)*
g3097 not 2743GAT(888) ; 2743GAT(888)*
g3098 not 2744GAT(889) ; 2744GAT(889)*
g3099 not 2739GAT(890) ; 2739GAT(890)*
g3100 not 2736GAT(891) ; 2736GAT(891)*
g3101 not 2733GAT(892) ; 2733GAT(892)*
g3102 not 2731GAT(893) ; 2731GAT(893)*
g3103 not 2732GAT(897) ; 2732GAT(897)*
g3104 not 2727GAT(899) ; 2727GAT(899)*
g3105 not 2724GAT(894) ; 2724GAT(894)*
g3106 not 1038GAT(122) ; 1038GAT(122)*
g3107 not 2721GAT(895) ; 2721GAT(895)*
g3108 not 990GAT(138) ; 990GAT(138)*
g3109 not 2718GAT(896) ; 2718GAT(896)*
g3110 not 942GAT(154) ; 942GAT(154)*
g3111 not 2715GAT(898) ; 2715GAT(898)*
g3112 not 894GAT(170) ; 894GAT(170)*
g3113 not 2712GAT(900) ; 2712GAT(900)*
g3114 not 846GAT(186) ; 846GAT(186)*
g3115 not 2709GAT(901) ; 2709GAT(901)*
g3116 not 798GAT(202) ; 798GAT(202)*
g3117 not 2706GAT(902) ; 2706GAT(902)*
g3118 not 750GAT(218) ; 750GAT(218)*
g3119 not 2703GAT(903) ; 2703GAT(903)*
g3120 not 702GAT(234) ; 702GAT(234)*
g3121 not 2700GAT(904) ; 2700GAT(904)*
g3122 not 654GAT(250) ; 654GAT(250)*
g3123 not 2697GAT(905) ; 2697GAT(905)*
g3124 not 606GAT(266) ; 606GAT(266)*
g3125 not 2694GAT(906) ; 2694GAT(906)*
g3126 not 558GAT(282) ; 558GAT(282)*
g3127 not 2801GAT(908) ; 2801GAT(908)*
g3128 not 2802GAT(909) ; 2802GAT(909)*
g3129 not 2797GAT(910) ; 2797GAT(910)*
g3130 not 2794GAT(911) ; 2794GAT(911)*
g3131 not 2791GAT(912) ; 2791GAT(912)*
g3132 not 2789GAT(913) ; 2789GAT(913)*
g3133 not 2790GAT(914) ; 2790GAT(914)*
g3134 not 2785GAT(915) ; 2785GAT(915)*
g3135 not 2803GAT(907) ; 2803GAT(907)*
g3136 not 1233GAT(57) ; 1233GAT(57)*
g3137 not 2781GAT(916) ; 2781GAT(916)*
g3138 not 2777GAT(917) ; 2777GAT(917)*
g3139 not 2773GAT(918) ; 2773GAT(918)*
g3140 not 2769GAT(919) ; 2769GAT(919)*
g3141 not 2765GAT(920) ; 2765GAT(920)*
g3142 not 2761GAT(921) ; 2761GAT(921)*
g3143 not 2757GAT(922) ; 2757GAT(922)*
g3144 not 2753GAT(923) ; 2753GAT(923)*
g3145 not 2749GAT(924) ; 2749GAT(924)*
g3146 not 2745GAT(925) ; 2745GAT(925)*
g3147 not 2873GAT(932) ; 2873GAT(932)*
g3148 not 2868GAT(927) ; 2868GAT(927)*
g3149 not 2869GAT(928) ; 2869GAT(928)*
g3150 not 2864GAT(929) ; 2864GAT(929)*
g3151 not 2861GAT(930) ; 2861GAT(930)*
g3152 not 2858GAT(936) ; 2858GAT(936)*
g3153 not 2856GAT(931) ; 2856GAT(931)*
g3154 not 2857GAT(938) ; 2857GAT(938)*
g3155 not 2851GAT(933) ; 2851GAT(933)*
g3156 not 2852GAT(941) ; 2852GAT(941)*
g3157 not 2870GAT(926) ; 2870GAT(926)*
g3158 not 1185GAT(73) ; 1185GAT(73)*
g3159 not 2846GAT(934) ; 2846GAT(934)*
g3160 not 2847GAT(944) ; 2847GAT(944)*
g3161 not 2841GAT(935) ; 2841GAT(935)*
g3162 not 2842GAT(947) ; 2842GAT(947)*
g3163 not 2836GAT(937) ; 2836GAT(937)*
g3164 not 2837GAT(950) ; 2837GAT(950)*
g3165 not 2831GAT(940) ; 2831GAT(940)*
g3166 not 2832GAT(953) ; 2832GAT(953)*
g3167 not 2826GAT(943) ; 2826GAT(943)*
g3168 not 2827GAT(956) ; 2827GAT(956)*
g3169 not 2821GAT(946) ; 2821GAT(946)*
g3170 not 2822GAT(958) ; 2822GAT(958)*
g3171 not 2816GAT(949) ; 2816GAT(949)*
g3172 not 2817GAT(960) ; 2817GAT(960)*
g3173 not 2811GAT(952) ; 2811GAT(952)*
g3174 not 2812GAT(962) ; 2812GAT(962)*
g3175 not 2806GAT(955) ; 2806GAT(955)*
g3176 not 2807GAT(964) ; 2807GAT(964)*
g3177 not 1281GAT(41) ; 1281GAT(41)*
g3178 not 2923GAT(965) ; 2923GAT(965)*
g3179 not 2921GAT(966) ; 2921GAT(966)*
g3180 not 2922GAT(972) ; 2922GAT(972)*
g3181 not 2917GAT(974) ; 2917GAT(974)*
g3182 not 2912GAT(968) ; 2912GAT(968)*
g3183 not 2913GAT(969) ; 2913GAT(969)*
g3184 not 2908GAT(970) ; 2908GAT(970)*
g3185 not 2914GAT(967) ; 2914GAT(967)*
g3186 not 1137GAT(89) ; 1137GAT(89)*
g3187 not 2905GAT(971) ; 2905GAT(971)*
g3188 not 2853GAT(939) ; 2853GAT(939)*
g3189 not 2902GAT(973) ; 2902GAT(973)*
g3190 not 2848GAT(942) ; 2848GAT(942)*
g3191 not 2899GAT(975) ; 2899GAT(975)*
g3192 not 2843GAT(945) ; 2843GAT(945)*
g3193 not 2896GAT(976) ; 2896GAT(976)*
g3194 not 2838GAT(948) ; 2838GAT(948)*
g3195 not 2893GAT(977) ; 2893GAT(977)*
g3196 not 2833GAT(951) ; 2833GAT(951)*
g3197 not 2890GAT(978) ; 2890GAT(978)*
g3198 not 2828GAT(954) ; 2828GAT(954)*
g3199 not 2887GAT(979) ; 2887GAT(979)*
g3200 not 2823GAT(957) ; 2823GAT(957)*
g3201 not 2884GAT(980) ; 2884GAT(980)*
g3202 not 2818GAT(959) ; 2818GAT(959)*
g3203 not 2881GAT(981) ; 2881GAT(981)*
g3204 not 2813GAT(961) ; 2813GAT(961)*
g3205 not 2878GAT(982) ; 2878GAT(982)*
g3206 not 2808GAT(963) ; 2808GAT(963)*
g3207 not 2983GAT(984) ; 2983GAT(984)*
g3208 not 2980GAT(985) ; 2980GAT(985)*
g3209 not 2977GAT(986) ; 2977GAT(986)*
g3210 not 2975GAT(987) ; 2975GAT(987)*
g3211 not 2976GAT(990) ; 2976GAT(990)*
g3212 not 2971GAT(991) ; 2971GAT(991)*
g3213 not 2966GAT(989) ; 2966GAT(989)*
g3214 not 2967GAT(992) ; 2967GAT(992)*
g3215 not 2962GAT(993) ; 2962GAT(993)*
g3216 not 2958GAT(994) ; 2958GAT(994)*
g3217 not 2954GAT(995) ; 2954GAT(995)*
g3218 not 2950GAT(996) ; 2950GAT(996)*
g3219 not 2968GAT(988) ; 2968GAT(988)*
g3220 not 1089GAT(105) ; 1089GAT(105)*
g3221 not 2946GAT(997) ; 2946GAT(997)*
g3222 not 2942GAT(998) ; 2942GAT(998)*
g3223 not 2938GAT(999) ; 2938GAT(999)*
g3224 not 2934GAT(1000) ; 2934GAT(1000)*
g3225 not 2930GAT(1001) ; 2930GAT(1001)*
g3226 not 2926GAT(1002) ; 2926GAT(1002)*
g3227 not 3026GAT(1003) ; 3026GAT(1003)*
g3228 not 3027GAT(1004) ; 3027GAT(1004)*
g3229 not 3022GAT(1005) ; 3022GAT(1005)*
g3230 not 3019GAT(1006) ; 3019GAT(1006)*
g3231 not 3016GAT(1007) ; 3016GAT(1007)*
g3232 not 3014GAT(1008) ; 3014GAT(1008)*
g3233 not 3015GAT(1013) ; 3015GAT(1013)*
g3234 not 3010GAT(1015) ; 3010GAT(1015)*
g3235 not 3005GAT(1010) ; 3005GAT(1010)*
g3236 not 3006GAT(1017) ; 3006GAT(1017)*
g3237 not 3003GAT(1011) ; 3003GAT(1011)*
g3238 not 3004GAT(1019) ; 3004GAT(1019)*
g3239 not 3001GAT(1012) ; 3001GAT(1012)*
g3240 not 3002GAT(1021) ; 3002GAT(1021)*
g3241 not 2999GAT(1014) ; 2999GAT(1014)*
g3242 not 3000GAT(1023) ; 3000GAT(1023)*
g3243 not 2997GAT(1016) ; 2997GAT(1016)*
g3244 not 2998GAT(1025) ; 2998GAT(1025)*
g3245 not 3007GAT(1009) ; 3007GAT(1009)*
g3246 not 1041GAT(121) ; 1041GAT(121)*
g3247 not 2995GAT(1018) ; 2995GAT(1018)*
g3248 not 2996GAT(1027) ; 2996GAT(1027)*
g3249 not 2993GAT(1020) ; 2993GAT(1020)*
g3250 not 2994GAT(1028) ; 2994GAT(1028)*
g3251 not 2991GAT(1022) ; 2991GAT(1022)*
g3252 not 2992GAT(1029) ; 2992GAT(1029)*
g3253 not 2989GAT(1024) ; 2989GAT(1024)*
g3254 not 2990GAT(1030) ; 2990GAT(1030)*
g3255 not 2987GAT(1026) ; 2987GAT(1026)*
g3256 not 2988GAT(1031) ; 2988GAT(1031)*
g3257 not 3074GAT(1033) ; 3074GAT(1033)*
g3258 not 3075GAT(1034) ; 3075GAT(1034)*
g3259 not 3070GAT(1035) ; 3070GAT(1035)*
g3260 not 3067GAT(1036) ; 3067GAT(1036)*
g3261 not 3064GAT(1037) ; 3064GAT(1037)*
g3262 not 3062GAT(1038) ; 3062GAT(1038)*
g3263 not 3063GAT(1043) ; 3063GAT(1043)*
g3264 not 3058GAT(1045) ; 3058GAT(1045)*
g3265 not 3076GAT(1032) ; 3076GAT(1032)*
g3266 not 1236GAT(56) ; 1236GAT(56)*
g3267 not 3055GAT(1039) ; 3055GAT(1039)*
g3268 not 993GAT(137) ; 993GAT(137)*
g3269 not 3052GAT(1040) ; 3052GAT(1040)*
g3270 not 945GAT(153) ; 945GAT(153)*
g3271 not 3049GAT(1041) ; 3049GAT(1041)*
g3272 not 897GAT(169) ; 897GAT(169)*
g3273 not 3046GAT(1042) ; 3046GAT(1042)*
g3274 not 849GAT(185) ; 849GAT(185)*
g3275 not 3043GAT(1044) ; 3043GAT(1044)*
g3276 not 801GAT(201) ; 801GAT(201)*
g3277 not 3040GAT(1046) ; 3040GAT(1046)*
g3278 not 753GAT(217) ; 753GAT(217)*
g3279 not 3037GAT(1047) ; 3037GAT(1047)*
g3280 not 705GAT(233) ; 705GAT(233)*
g3281 not 3034GAT(1048) ; 3034GAT(1048)*
g3282 not 657GAT(249) ; 657GAT(249)*
g3283 not 3031GAT(1049) ; 3031GAT(1049)*
g3284 not 609GAT(265) ; 609GAT(265)*
g3285 not 3028GAT(1050) ; 3028GAT(1050)*
g3286 not 561GAT(281) ; 561GAT(281)*
g3287 not 3136GAT(1058) ; 3136GAT(1058)*
g3288 not 3131GAT(1052) ; 3131GAT(1052)*
g3289 not 3132GAT(1053) ; 3132GAT(1053)*
g3290 not 3127GAT(1054) ; 3127GAT(1054)*
g3291 not 3124GAT(1055) ; 3124GAT(1055)*
g3292 not 3121GAT(1056) ; 3121GAT(1056)*
g3293 not 3119GAT(1057) ; 3119GAT(1057)*
g3294 not 3120GAT(1059) ; 3120GAT(1059)*
g3295 not 3115GAT(1060) ; 3115GAT(1060)*
g3296 not 3111GAT(1061) ; 3111GAT(1061)*
g3297 not 3133GAT(1051) ; 3133GAT(1051)*
g3298 not 1188GAT(72) ; 1188GAT(72)*
g3299 not 3107GAT(1062) ; 3107GAT(1062)*
g3300 not 3103GAT(1063) ; 3103GAT(1063)*
g3301 not 3099GAT(1064) ; 3099GAT(1064)*
g3302 not 3095GAT(1065) ; 3095GAT(1065)*
g3303 not 3091GAT(1066) ; 3091GAT(1066)*
g3304 not 3087GAT(1067) ; 3087GAT(1067)*
g3305 not 3083GAT(1068) ; 3083GAT(1068)*
g3306 not 3079GAT(1069) ; 3079GAT(1069)*
g3307 not 1284GAT(40) ; 1284GAT(40)*
g3308 not 3208GAT(1070) ; 3208GAT(1070)*
g3309 not 3206GAT(1071) ; 3206GAT(1071)*
g3310 not 3207GAT(1078) ; 3207GAT(1078)*
g3311 not 3202GAT(1080) ; 3202GAT(1080)*
g3312 not 3197GAT(1073) ; 3197GAT(1073)*
g3313 not 3198GAT(1074) ; 3198GAT(1074)*
g3314 not 3193GAT(1075) ; 3193GAT(1075)*
g3315 not 3190GAT(1076) ; 3190GAT(1076)*
g3316 not 3187GAT(1084) ; 3187GAT(1084)*
g3317 not 3185GAT(1077) ; 3185GAT(1077)*
g3318 not 3186GAT(1086) ; 3186GAT(1086)*
g3319 not 3180GAT(1079) ; 3180GAT(1079)*
g3320 not 3181GAT(1089) ; 3181GAT(1089)*
g3321 not 3175GAT(1081) ; 3175GAT(1081)*
g3322 not 3176GAT(1092) ; 3176GAT(1092)*
g3323 not 3199GAT(1072) ; 3199GAT(1072)*
g3324 not 1140GAT(88) ; 1140GAT(88)*
g3325 not 3170GAT(1082) ; 3170GAT(1082)*
g3326 not 3171GAT(1095) ; 3171GAT(1095)*
g3327 not 3165GAT(1083) ; 3165GAT(1083)*
g3328 not 3166GAT(1098) ; 3166GAT(1098)*
g3329 not 3160GAT(1085) ; 3160GAT(1085)*
g3330 not 3161GAT(1100) ; 3161GAT(1100)*
g3331 not 3155GAT(1088) ; 3155GAT(1088)*
g3332 not 3156GAT(1102) ; 3156GAT(1102)*
g3333 not 3150GAT(1091) ; 3150GAT(1091)*
g3334 not 3151GAT(1104) ; 3151GAT(1104)*
g3335 not 3145GAT(1094) ; 3145GAT(1094)*
g3336 not 3146GAT(1106) ; 3146GAT(1106)*
g3337 not 3140GAT(1097) ; 3140GAT(1097)*
g3338 not 3141GAT(1108) ; 3141GAT(1108)*
g3339 not 3260GAT(1109) ; 3260GAT(1109)*
g3340 not 3257GAT(1110) ; 3257GAT(1110)*
g3341 not 3254GAT(1111) ; 3254GAT(1111)*
g3342 not 3252GAT(1112) ; 3252GAT(1112)*
g3343 not 3253GAT(1119) ; 3253GAT(1119)*
g3344 not 3248GAT(1121) ; 3248GAT(1121)*
g3345 not 3243GAT(1114) ; 3243GAT(1114)*
g3346 not 3244GAT(1115) ; 3244GAT(1115)*
g3347 not 3239GAT(1116) ; 3239GAT(1116)*
g3348 not 3245GAT(1113) ; 3245GAT(1113)*
g3349 not 1092GAT(104) ; 1092GAT(104)*
g3350 not 3236GAT(1117) ; 3236GAT(1117)*
g3351 not 3182GAT(1087) ; 3182GAT(1087)*
g3352 not 3233GAT(1118) ; 3233GAT(1118)*
g3353 not 3177GAT(1090) ; 3177GAT(1090)*
g3354 not 3230GAT(1120) ; 3230GAT(1120)*
g3355 not 3172GAT(1093) ; 3172GAT(1093)*
g3356 not 3227GAT(1122) ; 3227GAT(1122)*
g3357 not 3167GAT(1096) ; 3167GAT(1096)*
g3358 not 3224GAT(1123) ; 3224GAT(1123)*
g3359 not 3162GAT(1099) ; 3162GAT(1099)*
g3360 not 3221GAT(1124) ; 3221GAT(1124)*
g3361 not 3157GAT(1101) ; 3157GAT(1101)*
g3362 not 3218GAT(1125) ; 3218GAT(1125)*
g3363 not 3152GAT(1103) ; 3152GAT(1103)*
g3364 not 3215GAT(1126) ; 3215GAT(1126)*
g3365 not 3147GAT(1105) ; 3147GAT(1105)*
g3366 not 3212GAT(1127) ; 3212GAT(1127)*
g3367 not 3142GAT(1107) ; 3142GAT(1107)*
g3368 not 3321GAT(1129) ; 3321GAT(1129)*
g3369 not 3322GAT(1130) ; 3322GAT(1130)*
g3370 not 3317GAT(1131) ; 3317GAT(1131)*
g3371 not 3314GAT(1132) ; 3314GAT(1132)*
g3372 not 3311GAT(1133) ; 3311GAT(1133)*
g3373 not 3309GAT(1134) ; 3309GAT(1134)*
g3374 not 3310GAT(1137) ; 3310GAT(1137)*
g3375 not 3305GAT(1138) ; 3305GAT(1138)*
g3376 not 3300GAT(1136) ; 3300GAT(1136)*
g3377 not 3301GAT(1139) ; 3301GAT(1139)*
g3378 not 3296GAT(1140) ; 3296GAT(1140)*
g3379 not 3292GAT(1141) ; 3292GAT(1141)*
g3380 not 3288GAT(1142) ; 3288GAT(1142)*
g3381 not 3284GAT(1143) ; 3284GAT(1143)*
g3382 not 3280GAT(1144) ; 3280GAT(1144)*
g3383 not 3302GAT(1135) ; 3302GAT(1135)*
g3384 not 1044GAT(120) ; 1044GAT(120)*
g3385 not 3276GAT(1145) ; 3276GAT(1145)*
g3386 not 3272GAT(1146) ; 3272GAT(1146)*
g3387 not 3268GAT(1147) ; 3268GAT(1147)*
g3388 not 3264GAT(1148) ; 3264GAT(1148)*
g3389 not 3360GAT(1150) ; 3360GAT(1150)*
g3390 not 3361GAT(1151) ; 3361GAT(1151)*
g3391 not 3356GAT(1152) ; 3356GAT(1152)*
g3392 not 3353GAT(1153) ; 3353GAT(1153)*
g3393 not 3350GAT(1154) ; 3350GAT(1154)*
g3394 not 3348GAT(1155) ; 3348GAT(1155)*
g3395 not 3349GAT(1161) ; 3349GAT(1161)*
g3396 not 3344GAT(1163) ; 3344GAT(1163)*
g3397 not 3339GAT(1157) ; 3339GAT(1157)*
g3398 not 3340GAT(1165) ; 3340GAT(1165)*
g3399 not 3362GAT(1149) ; 3362GAT(1149)*
g3400 not 1239GAT(55) ; 1239GAT(55)*
g3401 not 3337GAT(1158) ; 3337GAT(1158)*
g3402 not 3338GAT(1167) ; 3338GAT(1167)*
g3403 not 3335GAT(1159) ; 3335GAT(1159)*
g3404 not 3336GAT(1169) ; 3336GAT(1169)*
g3405 not 3333GAT(1160) ; 3333GAT(1160)*
g3406 not 3334GAT(1171) ; 3334GAT(1171)*
g3407 not 3331GAT(1162) ; 3331GAT(1162)*
g3408 not 3332GAT(1172) ; 3332GAT(1172)*
g3409 not 3329GAT(1164) ; 3329GAT(1164)*
g3410 not 3330GAT(1173) ; 3330GAT(1173)*
g3411 not 3341GAT(1156) ; 3341GAT(1156)*
g3412 not 996GAT(136) ; 996GAT(136)*
g3413 not 3327GAT(1166) ; 3327GAT(1166)*
g3414 not 3328GAT(1174) ; 3328GAT(1174)*
g3415 not 3325GAT(1168) ; 3325GAT(1168)*
g3416 not 3326GAT(1175) ; 3326GAT(1175)*
g3417 not 3323GAT(1170) ; 3323GAT(1170)*
g3418 not 3324GAT(1176) ; 3324GAT(1176)*
g3419 not 3413GAT(1185) ; 3413GAT(1185)*
g3420 not 3408GAT(1178) ; 3408GAT(1178)*
g3421 not 3409GAT(1179) ; 3409GAT(1179)*
g3422 not 3404GAT(1180) ; 3404GAT(1180)*
g3423 not 3401GAT(1181) ; 3401GAT(1181)*
g3424 not 3398GAT(1182) ; 3398GAT(1182)*
g3425 not 3396GAT(1183) ; 3396GAT(1183)*
g3426 not 3397GAT(1190) ; 3397GAT(1190)*
g3427 not 3392GAT(1192) ; 3392GAT(1192)*
g3428 not 3410GAT(1177) ; 3410GAT(1177)*
g3429 not 1191GAT(71) ; 1191GAT(71)*
g3430 not 3389GAT(1184) ; 3389GAT(1184)*
g3431 not 948GAT(152) ; 948GAT(152)*
g3432 not 3386GAT(1186) ; 3386GAT(1186)*
g3433 not 900GAT(168) ; 900GAT(168)*
g3434 not 3383GAT(1187) ; 3383GAT(1187)*
g3435 not 852GAT(184) ; 852GAT(184)*
g3436 not 3380GAT(1188) ; 3380GAT(1188)*
g3437 not 804GAT(200) ; 804GAT(200)*
g3438 not 3377GAT(1189) ; 3377GAT(1189)*
g3439 not 756GAT(216) ; 756GAT(216)*
g3440 not 3374GAT(1191) ; 3374GAT(1191)*
g3441 not 708GAT(232) ; 708GAT(232)*
g3442 not 3371GAT(1193) ; 3371GAT(1193)*
g3443 not 660GAT(248) ; 660GAT(248)*
g3444 not 3368GAT(1194) ; 3368GAT(1194)*
g3445 not 612GAT(264) ; 612GAT(264)*
g3446 not 3365GAT(1195) ; 3365GAT(1195)*
g3447 not 564GAT(280) ; 564GAT(280)*
g3448 not 1287GAT(39) ; 1287GAT(39)*
g3449 not 3476GAT(1196) ; 3476GAT(1196)*
g3450 not 3474GAT(1197) ; 3474GAT(1197)*
g3451 not 3475GAT(1205) ; 3475GAT(1205)*
g3452 not 3470GAT(1206) ; 3470GAT(1206)*
g3453 not 3465GAT(1199) ; 3465GAT(1199)*
g3454 not 3466GAT(1200) ; 3466GAT(1200)*
g3455 not 3461GAT(1201) ; 3461GAT(1201)*
g3456 not 3458GAT(1202) ; 3458GAT(1202)*
g3457 not 3455GAT(1203) ; 3455GAT(1203)*
g3458 not 3453GAT(1204) ; 3453GAT(1204)*
g3459 not 3454GAT(1207) ; 3454GAT(1207)*
g3460 not 3449GAT(1208) ; 3449GAT(1208)*
g3461 not 3445GAT(1209) ; 3445GAT(1209)*
g3462 not 3441GAT(1210) ; 3441GAT(1210)*
g3463 not 3467GAT(1198) ; 3467GAT(1198)*
g3464 not 1143GAT(87) ; 1143GAT(87)*
g3465 not 3437GAT(1211) ; 3437GAT(1211)*
g3466 not 3433GAT(1212) ; 3433GAT(1212)*
g3467 not 3429GAT(1213) ; 3429GAT(1213)*
g3468 not 3425GAT(1214) ; 3425GAT(1214)*
g3469 not 3421GAT(1215) ; 3421GAT(1215)*
g3470 not 3417GAT(1216) ; 3417GAT(1216)*
g3471 not 3548GAT(1217) ; 3548GAT(1217)*
g3472 not 3545GAT(1218) ; 3545GAT(1218)*
g3473 not 3542GAT(1219) ; 3542GAT(1219)*
g3474 not 3540GAT(1220) ; 3540GAT(1220)*
g3475 not 3541GAT(1228) ; 3541GAT(1228)*
g3476 not 3536GAT(1230) ; 3536GAT(1230)*
g3477 not 3531GAT(1222) ; 3531GAT(1222)*
g3478 not 3532GAT(1223) ; 3532GAT(1223)*
g3479 not 3527GAT(1224) ; 3527GAT(1224)*
g3480 not 3524GAT(1225) ; 3524GAT(1225)*
g3481 not 3521GAT(1234) ; 3521GAT(1234)*
g3482 not 3519GAT(1226) ; 3519GAT(1226)*
g3483 not 3520GAT(1236) ; 3520GAT(1236)*
g3484 not 3514GAT(1227) ; 3514GAT(1227)*
g3485 not 3515GAT(1239) ; 3515GAT(1239)*
g3486 not 3509GAT(1229) ; 3509GAT(1229)*
g3487 not 3510GAT(1242) ; 3510GAT(1242)*
g3488 not 3504GAT(1231) ; 3504GAT(1231)*
g3489 not 3505GAT(1244) ; 3505GAT(1244)*
g3490 not 3533GAT(1221) ; 3533GAT(1221)*
g3491 not 1095GAT(103) ; 1095GAT(103)*
g3492 not 3499GAT(1232) ; 3499GAT(1232)*
g3493 not 3500GAT(1246) ; 3500GAT(1246)*
g3494 not 3494GAT(1233) ; 3494GAT(1233)*
g3495 not 3495GAT(1248) ; 3495GAT(1248)*
g3496 not 3489GAT(1235) ; 3489GAT(1235)*
g3497 not 3490GAT(1250) ; 3490GAT(1250)*
g3498 not 3484GAT(1238) ; 3484GAT(1238)*
g3499 not 3485GAT(1252) ; 3485GAT(1252)*
g3500 not 3479GAT(1241) ; 3479GAT(1241)*
g3501 not 3480GAT(1254) ; 3480GAT(1254)*
g3502 not 3602GAT(1255) ; 3602GAT(1255)*
g3503 not 3603GAT(1256) ; 3603GAT(1256)*
g3504 not 3598GAT(1257) ; 3598GAT(1257)*
g3505 not 3595GAT(1258) ; 3595GAT(1258)*
g3506 not 3592GAT(1259) ; 3592GAT(1259)*
g3507 not 3590GAT(1260) ; 3590GAT(1260)*
g3508 not 3591GAT(1268) ; 3591GAT(1268)*
g3509 not 3586GAT(1270) ; 3586GAT(1270)*
g3510 not 3581GAT(1262) ; 3581GAT(1262)*
g3511 not 3582GAT(1263) ; 3582GAT(1263)*
g3512 not 3577GAT(1264) ; 3577GAT(1264)*
g3513 not 3583GAT(1261) ; 3583GAT(1261)*
g3514 not 1047GAT(119) ; 1047GAT(119)*
g3515 not 3574GAT(1265) ; 3574GAT(1265)*
g3516 not 3516GAT(1237) ; 3516GAT(1237)*
g3517 not 3571GAT(1266) ; 3571GAT(1266)*
g3518 not 3511GAT(1240) ; 3511GAT(1240)*
g3519 not 3568GAT(1267) ; 3568GAT(1267)*
g3520 not 3506GAT(1243) ; 3506GAT(1243)*
g3521 not 3565GAT(1269) ; 3565GAT(1269)*
g3522 not 3501GAT(1245) ; 3501GAT(1245)*
g3523 not 3562GAT(1271) ; 3562GAT(1271)*
g3524 not 3496GAT(1247) ; 3496GAT(1247)*
g3525 not 3559GAT(1272) ; 3559GAT(1272)*
g3526 not 3491GAT(1249) ; 3491GAT(1249)*
g3527 not 3556GAT(1273) ; 3556GAT(1273)*
g3528 not 3486GAT(1251) ; 3486GAT(1251)*
g3529 not 3553GAT(1274) ; 3553GAT(1274)*
g3530 not 3481GAT(1253) ; 3481GAT(1253)*
g3531 not 3657GAT(1277) ; 3657GAT(1277)*
g3532 not 3658GAT(1278) ; 3658GAT(1278)*
g3533 not 3653GAT(1279) ; 3653GAT(1279)*
g3534 not 3650GAT(1280) ; 3650GAT(1280)*
g3535 not 3647GAT(1281) ; 3647GAT(1281)*
g3536 not 3645GAT(1282) ; 3645GAT(1282)*
g3537 not 3646GAT(1285) ; 3646GAT(1285)*
g3538 not 3641GAT(1286) ; 3641GAT(1286)*
g3539 not 3636GAT(1284) ; 3636GAT(1284)*
g3540 not 3637GAT(1287) ; 3637GAT(1287)*
g3541 not 3632GAT(1288) ; 3632GAT(1288)*
g3542 not 3659GAT(1276) ; 3659GAT(1276)*
g3543 not 1242GAT(54) ; 1242GAT(54)*
g3544 not 3628GAT(1289) ; 3628GAT(1289)*
g3545 not 3624GAT(1290) ; 3624GAT(1290)*
g3546 not 3620GAT(1291) ; 3620GAT(1291)*
g3547 not 3616GAT(1292) ; 3616GAT(1292)*
g3548 not 3612GAT(1293) ; 3612GAT(1293)*
g3549 not 3638GAT(1283) ; 3638GAT(1283)*
g3550 not 999GAT(135) ; 999GAT(135)*
g3551 not 3608GAT(1294) ; 3608GAT(1294)*
g3552 not 3604GAT(1295) ; 3604GAT(1295)*
g3553 not 3702GAT(1305) ; 3702GAT(1305)*
g3554 not 3697GAT(1297) ; 3697GAT(1297)*
g3555 not 3698GAT(1298) ; 3698GAT(1298)*
g3556 not 3693GAT(1299) ; 3693GAT(1299)*
g3557 not 3690GAT(1300) ; 3690GAT(1300)*
g3558 not 3687GAT(1301) ; 3687GAT(1301)*
g3559 not 3685GAT(1302) ; 3685GAT(1302)*
g3560 not 3686GAT(1310) ; 3686GAT(1310)*
g3561 not 3681GAT(1312) ; 3681GAT(1312)*
g3562 not 3676GAT(1304) ; 3676GAT(1304)*
g3563 not 3677GAT(1314) ; 3677GAT(1314)*
g3564 not 3674GAT(1306) ; 3674GAT(1306)*
g3565 not 3675GAT(1316) ; 3675GAT(1316)*
g3566 not 3699GAT(1296) ; 3699GAT(1296)*
g3567 not 1194GAT(70) ; 1194GAT(70)*
g3568 not 3672GAT(1307) ; 3672GAT(1307)*
g3569 not 3673GAT(1317) ; 3673GAT(1317)*
g3570 not 3670GAT(1308) ; 3670GAT(1308)*
g3571 not 3671GAT(1318) ; 3671GAT(1318)*
g3572 not 3668GAT(1309) ; 3668GAT(1309)*
g3573 not 3669GAT(1319) ; 3669GAT(1319)*
g3574 not 3666GAT(1311) ; 3666GAT(1311)*
g3575 not 3667GAT(1320) ; 3667GAT(1320)*
g3576 not 3664GAT(1313) ; 3664GAT(1313)*
g3577 not 3665GAT(1321) ; 3665GAT(1321)*
g3578 not 3678GAT(1303) ; 3678GAT(1303)*
g3579 not 951GAT(151) ; 951GAT(151)*
g3580 not 3662GAT(1315) ; 3662GAT(1315)*
g3581 not 3663GAT(1322) ; 3663GAT(1322)*
g3582 not 1290GAT(38) ; 1290GAT(38)*
g3583 not 3757GAT(1323) ; 3757GAT(1323)*
g3584 not 3755GAT(1324) ; 3755GAT(1324)*
g3585 not 3756GAT(1333) ; 3756GAT(1333)*
g3586 not 3751GAT(1335) ; 3751GAT(1335)*
g3587 not 3746GAT(1326) ; 3746GAT(1326)*
g3588 not 3747GAT(1327) ; 3747GAT(1327)*
g3589 not 3742GAT(1328) ; 3742GAT(1328)*
g3590 not 3739GAT(1329) ; 3739GAT(1329)*
g3591 not 3736GAT(1330) ; 3736GAT(1330)*
g3592 not 3734GAT(1331) ; 3734GAT(1331)*
g3593 not 3735GAT(1340) ; 3735GAT(1340)*
g3594 not 3730GAT(1342) ; 3730GAT(1342)*
g3595 not 3748GAT(1325) ; 3748GAT(1325)*
g3596 not 1146GAT(86) ; 1146GAT(86)*
g3597 not 3727GAT(1332) ; 3727GAT(1332)*
g3598 not 903GAT(167) ; 903GAT(167)*
g3599 not 3724GAT(1334) ; 3724GAT(1334)*
g3600 not 855GAT(183) ; 855GAT(183)*
g3601 not 3721GAT(1336) ; 3721GAT(1336)*
g3602 not 807GAT(199) ; 807GAT(199)*
g3603 not 3718GAT(1337) ; 3718GAT(1337)*
g3604 not 759GAT(215) ; 759GAT(215)*
g3605 not 3715GAT(1338) ; 3715GAT(1338)*
g3606 not 711GAT(231) ; 711GAT(231)*
g3607 not 3712GAT(1339) ; 3712GAT(1339)*
g3608 not 663GAT(247) ; 663GAT(247)*
g3609 not 3709GAT(1341) ; 3709GAT(1341)*
g3610 not 615GAT(263) ; 615GAT(263)*
g3611 not 3706GAT(1343) ; 3706GAT(1343)*
g3612 not 567GAT(279) ; 567GAT(279)*
g3613 not 3821GAT(1344) ; 3821GAT(1344)*
g3614 not 3818GAT(1345) ; 3818GAT(1345)*
g3615 not 3815GAT(1346) ; 3815GAT(1346)*
g3616 not 3813GAT(1347) ; 3813GAT(1347)*
g3617 not 3814GAT(1355) ; 3814GAT(1355)*
g3618 not 3809GAT(1356) ; 3809GAT(1356)*
g3619 not 3804GAT(1349) ; 3804GAT(1349)*
g3620 not 3805GAT(1350) ; 3805GAT(1350)*
g3621 not 3800GAT(1351) ; 3800GAT(1351)*
g3622 not 3797GAT(1352) ; 3797GAT(1352)*
g3623 not 3794GAT(1353) ; 3794GAT(1353)*
g3624 not 3792GAT(1354) ; 3792GAT(1354)*
g3625 not 3793GAT(1357) ; 3793GAT(1357)*
g3626 not 3788GAT(1358) ; 3788GAT(1358)*
g3627 not 3784GAT(1359) ; 3784GAT(1359)*
g3628 not 3780GAT(1360) ; 3780GAT(1360)*
g3629 not 3776GAT(1361) ; 3776GAT(1361)*
g3630 not 3806GAT(1348) ; 3806GAT(1348)*
g3631 not 1098GAT(102) ; 1098GAT(102)*
g3632 not 3772GAT(1362) ; 3772GAT(1362)*
g3633 not 3768GAT(1363) ; 3768GAT(1363)*
g3634 not 3764GAT(1364) ; 3764GAT(1364)*
g3635 not 3760GAT(1365) ; 3760GAT(1365)*
g3636 not 3893GAT(1366) ; 3893GAT(1366)*
g3637 not 3894GAT(1367) ; 3894GAT(1367)*
g3638 not 3889GAT(1368) ; 3889GAT(1368)*
g3639 not 3886GAT(1369) ; 3886GAT(1369)*
g3640 not 3883GAT(1370) ; 3883GAT(1370)*
g3641 not 3881GAT(1371) ; 3881GAT(1371)*
g3642 not 3882GAT(1380) ; 3882GAT(1380)*
g3643 not 3877GAT(1382) ; 3877GAT(1382)*
g3644 not 3872GAT(1373) ; 3872GAT(1373)*
g3645 not 3873GAT(1374) ; 3873GAT(1374)*
g3646 not 3868GAT(1375) ; 3868GAT(1375)*
g3647 not 3865GAT(1376) ; 3865GAT(1376)*
g3648 not 3862GAT(1386) ; 3862GAT(1386)*
g3649 not 3860GAT(1377) ; 3860GAT(1377)*
g3650 not 3861GAT(1388) ; 3861GAT(1388)*
g3651 not 3855GAT(1378) ; 3855GAT(1378)*
g3652 not 3856GAT(1390) ; 3856GAT(1390)*
g3653 not 3850GAT(1379) ; 3850GAT(1379)*
g3654 not 3851GAT(1392) ; 3851GAT(1392)*
g3655 not 3845GAT(1381) ; 3845GAT(1381)*
g3656 not 3846GAT(1394) ; 3846GAT(1394)*
g3657 not 3840GAT(1383) ; 3840GAT(1383)*
g3658 not 3841GAT(1396) ; 3841GAT(1396)*
g3659 not 3874GAT(1372) ; 3874GAT(1372)*
g3660 not 1050GAT(118) ; 1050GAT(118)*
g3661 not 3835GAT(1384) ; 3835GAT(1384)*
g3662 not 3836GAT(1398) ; 3836GAT(1398)*
g3663 not 3830GAT(1385) ; 3830GAT(1385)*
g3664 not 3831GAT(1400) ; 3831GAT(1400)*
g3665 not 3825GAT(1387) ; 3825GAT(1387)*
g3666 not 3826GAT(1402) ; 3826GAT(1402)*
g3667 not 3942GAT(1404) ; 3942GAT(1404)*
g3668 not 3943GAT(1405) ; 3943GAT(1405)*
g3669 not 3938GAT(1406) ; 3938GAT(1406)*
g3670 not 3935GAT(1407) ; 3935GAT(1407)*
g3671 not 3932GAT(1408) ; 3932GAT(1408)*
g3672 not 3930GAT(1409) ; 3930GAT(1409)*
g3673 not 3931GAT(1418) ; 3931GAT(1418)*
g3674 not 3926GAT(1420) ; 3926GAT(1420)*
g3675 not 3921GAT(1411) ; 3921GAT(1411)*
g3676 not 3922GAT(1412) ; 3922GAT(1412)*
g3677 not 3917GAT(1413) ; 3917GAT(1413)*
g3678 not 3944GAT(1403) ; 3944GAT(1403)*
g3679 not 1245GAT(53) ; 1245GAT(53)*
g3680 not 3923GAT(1410) ; 3923GAT(1410)*
g3681 not 1002GAT(134) ; 1002GAT(134)*
g3682 not 3914GAT(1414) ; 3914GAT(1414)*
g3683 not 3857GAT(1389) ; 3857GAT(1389)*
g3684 not 3911GAT(1415) ; 3911GAT(1415)*
g3685 not 3852GAT(1391) ; 3852GAT(1391)*
g3686 not 3908GAT(1416) ; 3908GAT(1416)*
g3687 not 3847GAT(1393) ; 3847GAT(1393)*
g3688 not 3905GAT(1417) ; 3905GAT(1417)*
g3689 not 3842GAT(1395) ; 3842GAT(1395)*
g3690 not 3902GAT(1419) ; 3902GAT(1419)*
g3691 not 3837GAT(1397) ; 3837GAT(1397)*
g3692 not 3899GAT(1421) ; 3899GAT(1421)*
g3693 not 3832GAT(1399) ; 3832GAT(1399)*
g3694 not 3896GAT(1422) ; 3896GAT(1422)*
g3695 not 3827GAT(1401) ; 3827GAT(1401)*
g3696 not 4001GAT(1433) ; 4001GAT(1433)*
g3697 not 3996GAT(1425) ; 3996GAT(1425)*
g3698 not 3997GAT(1426) ; 3997GAT(1426)*
g3699 not 3992GAT(1427) ; 3992GAT(1427)*
g3700 not 3989GAT(1428) ; 3989GAT(1428)*
g3701 not 3986GAT(1429) ; 3986GAT(1429)*
g3702 not 3984GAT(1430) ; 3984GAT(1430)*
g3703 not 3985GAT(1434) ; 3985GAT(1434)*
g3704 not 3980GAT(1435) ; 3980GAT(1435)*
g3705 not 3975GAT(1432) ; 3975GAT(1432)*
g3706 not 3976GAT(1436) ; 3976GAT(1436)*
g3707 not 3971GAT(1437) ; 3971GAT(1437)*
g3708 not 3967GAT(1438) ; 3967GAT(1438)*
g3709 not 3998GAT(1424) ; 3998GAT(1424)*
g3710 not 1197GAT(69) ; 1197GAT(69)*
g3711 not 3963GAT(1439) ; 3963GAT(1439)*
g3712 not 3959GAT(1440) ; 3959GAT(1440)*
g3713 not 3955GAT(1441) ; 3955GAT(1441)*
g3714 not 3951GAT(1442) ; 3951GAT(1442)*
g3715 not 3947GAT(1443) ; 3947GAT(1443)*
g3716 not 3977GAT(1431) ; 3977GAT(1431)*
g3717 not 954GAT(150) ; 954GAT(150)*
g3718 not 1293GAT(37) ; 1293GAT(37)*
g3719 not 4049GAT(1444) ; 4049GAT(1444)*
g3720 not 4047GAT(1445) ; 4047GAT(1445)*
g3721 not 4048GAT(1455) ; 4048GAT(1455)*
g3722 not 4043GAT(1457) ; 4043GAT(1457)*
g3723 not 4038GAT(1447) ; 4038GAT(1447)*
g3724 not 4039GAT(1448) ; 4039GAT(1448)*
g3725 not 4034GAT(1449) ; 4034GAT(1449)*
g3726 not 4031GAT(1450) ; 4031GAT(1450)*
g3727 not 4028GAT(1451) ; 4028GAT(1451)*
g3728 not 4026GAT(1452) ; 4026GAT(1452)*
g3729 not 4027GAT(1462) ; 4027GAT(1462)*
g3730 not 4022GAT(1464) ; 4022GAT(1464)*
g3731 not 4017GAT(1454) ; 4017GAT(1454)*
g3732 not 4018GAT(1465) ; 4018GAT(1465)*
g3733 not 4015GAT(1456) ; 4015GAT(1456)*
g3734 not 4016GAT(1466) ; 4016GAT(1466)*
g3735 not 4013GAT(1458) ; 4013GAT(1458)*
g3736 not 4014GAT(1467) ; 4014GAT(1467)*
g3737 not 4040GAT(1446) ; 4040GAT(1446)*
g3738 not 1149GAT(85) ; 1149GAT(85)*
g3739 not 4011GAT(1459) ; 4011GAT(1459)*
g3740 not 4012GAT(1468) ; 4012GAT(1468)*
g3741 not 4009GAT(1460) ; 4009GAT(1460)*
g3742 not 4010GAT(1469) ; 4010GAT(1469)*
g3743 not 4007GAT(1461) ; 4007GAT(1461)*
g3744 not 4008GAT(1470) ; 4008GAT(1470)*
g3745 not 4005GAT(1463) ; 4005GAT(1463)*
g3746 not 4006GAT(1471) ; 4006GAT(1471)*
g3747 not 4019GAT(1453) ; 4019GAT(1453)*
g3748 not 906GAT(166) ; 906GAT(166)*
g3749 not 4106GAT(1472) ; 4106GAT(1472)*
g3750 not 4103GAT(1473) ; 4103GAT(1473)*
g3751 not 4100GAT(1474) ; 4100GAT(1474)*
g3752 not 4098GAT(1475) ; 4098GAT(1475)*
g3753 not 4099GAT(1485) ; 4099GAT(1485)*
g3754 not 4094GAT(1487) ; 4094GAT(1487)*
g3755 not 4089GAT(1477) ; 4089GAT(1477)*
g3756 not 4090GAT(1478) ; 4090GAT(1478)*
g3757 not 4085GAT(1479) ; 4085GAT(1479)*
g3758 not 4082GAT(1480) ; 4082GAT(1480)*
g3759 not 4079GAT(1481) ; 4079GAT(1481)*
g3760 not 4077GAT(1482) ; 4077GAT(1482)*
g3761 not 4078GAT(1492) ; 4078GAT(1492)*
g3762 not 4073GAT(1493) ; 4073GAT(1493)*
g3763 not 4091GAT(1476) ; 4091GAT(1476)*
g3764 not 1101GAT(101) ; 1101GAT(101)*
g3765 not 4070GAT(1483) ; 4070GAT(1483)*
g3766 not 858GAT(182) ; 858GAT(182)*
g3767 not 4067GAT(1484) ; 4067GAT(1484)*
g3768 not 810GAT(198) ; 810GAT(198)*
g3769 not 4064GAT(1486) ; 4064GAT(1486)*
g3770 not 762GAT(214) ; 762GAT(214)*
g3771 not 4061GAT(1488) ; 4061GAT(1488)*
g3772 not 714GAT(230) ; 714GAT(230)*
g3773 not 4058GAT(1489) ; 4058GAT(1489)*
g3774 not 666GAT(246) ; 666GAT(246)*
g3775 not 4055GAT(1490) ; 4055GAT(1490)*
g3776 not 618GAT(262) ; 618GAT(262)*
g3777 not 4052GAT(1491) ; 4052GAT(1491)*
g3778 not 570GAT(278) ; 570GAT(278)*
g3779 not 4171GAT(1494) ; 4171GAT(1494)*
g3780 not 4172GAT(1495) ; 4172GAT(1495)*
g3781 not 4167GAT(1496) ; 4167GAT(1496)*
g3782 not 4164GAT(1497) ; 4164GAT(1497)*
g3783 not 4161GAT(1498) ; 4161GAT(1498)*
g3784 not 4159GAT(1499) ; 4159GAT(1499)*
g3785 not 4160GAT(1507) ; 4160GAT(1507)*
g3786 not 4155GAT(1508) ; 4155GAT(1508)*
g3787 not 4150GAT(1501) ; 4150GAT(1501)*
g3788 not 4151GAT(1502) ; 4151GAT(1502)*
g3789 not 4146GAT(1503) ; 4146GAT(1503)*
g3790 not 4143GAT(1504) ; 4143GAT(1504)*
g3791 not 4140GAT(1505) ; 4140GAT(1505)*
g3792 not 4138GAT(1506) ; 4138GAT(1506)*
g3793 not 4139GAT(1509) ; 4139GAT(1509)*
g3794 not 4134GAT(1510) ; 4134GAT(1510)*
g3795 not 4130GAT(1511) ; 4130GAT(1511)*
g3796 not 4126GAT(1512) ; 4126GAT(1512)*
g3797 not 4122GAT(1513) ; 4122GAT(1513)*
g3798 not 4118GAT(1514) ; 4118GAT(1514)*
g3799 not 4152GAT(1500) ; 4152GAT(1500)*
g3800 not 1053GAT(117) ; 1053GAT(117)*
g3801 not 4114GAT(1515) ; 4114GAT(1515)*
g3802 not 4110GAT(1516) ; 4110GAT(1516)*
g3803 not 4236GAT(1518) ; 4236GAT(1518)*
g3804 not 4237GAT(1519) ; 4237GAT(1519)*
g3805 not 4232GAT(1520) ; 4232GAT(1520)*
g3806 not 4229GAT(1521) ; 4229GAT(1521)*
g3807 not 4226GAT(1522) ; 4226GAT(1522)*
g3808 not 4224GAT(1523) ; 4224GAT(1523)*
g3809 not 4225GAT(1533) ; 4225GAT(1533)*
g3810 not 4220GAT(1535) ; 4220GAT(1535)*
g3811 not 4215GAT(1525) ; 4215GAT(1525)*
g3812 not 4216GAT(1526) ; 4216GAT(1526)*
g3813 not 4211GAT(1527) ; 4211GAT(1527)*
g3814 not 4208GAT(1528) ; 4208GAT(1528)*
g3815 not 4205GAT(1538) ; 4205GAT(1538)*
g3816 not 4203GAT(1529) ; 4203GAT(1529)*
g3817 not 4204GAT(1539) ; 4204GAT(1539)*
g3818 not 4238GAT(1517) ; 4238GAT(1517)*
g3819 not 1248GAT(52) ; 1248GAT(52)*
g3820 not 4198GAT(1530) ; 4198GAT(1530)*
g3821 not 4199GAT(1541) ; 4199GAT(1541)*
g3822 not 4193GAT(1531) ; 4193GAT(1531)*
g3823 not 4194GAT(1543) ; 4194GAT(1543)*
g3824 not 4188GAT(1532) ; 4188GAT(1532)*
g3825 not 4189GAT(1545) ; 4189GAT(1545)*
g3826 not 4183GAT(1534) ; 4183GAT(1534)*
g3827 not 4184GAT(1547) ; 4184GAT(1547)*
g3828 not 4178GAT(1536) ; 4178GAT(1536)*
g3829 not 4179GAT(1549) ; 4179GAT(1549)*
g3830 not 4217GAT(1524) ; 4217GAT(1524)*
g3831 not 1005GAT(133) ; 1005GAT(133)*
g3832 not 4173GAT(1537) ; 4173GAT(1537)*
g3833 not 4174GAT(1551) ; 4174GAT(1551)*
g3834 not 4290GAT(1564) ; 4290GAT(1564)*
g3835 not 4285GAT(1553) ; 4285GAT(1553)*
g3836 not 4286GAT(1554) ; 4286GAT(1554)*
g3837 not 4281GAT(1555) ; 4281GAT(1555)*
g3838 not 4278GAT(1556) ; 4278GAT(1556)*
g3839 not 4275GAT(1557) ; 4275GAT(1557)*
g3840 not 4273GAT(1558) ; 4273GAT(1558)*
g3841 not 4274GAT(1569) ; 4274GAT(1569)*
g3842 not 4269GAT(1571) ; 4269GAT(1571)*
g3843 not 4264GAT(1560) ; 4264GAT(1560)*
g3844 not 4265GAT(1561) ; 4265GAT(1561)*
g3845 not 4260GAT(1562) ; 4260GAT(1562)*
g3846 not 4287GAT(1552) ; 4287GAT(1552)*
g3847 not 1200GAT(68) ; 1200GAT(68)*
g3848 not 4266GAT(1559) ; 4266GAT(1559)*
g3849 not 957GAT(149) ; 957GAT(149)*
g3850 not 4257GAT(1563) ; 4257GAT(1563)*
g3851 not 4200GAT(1540) ; 4200GAT(1540)*
g3852 not 4254GAT(1565) ; 4254GAT(1565)*
g3853 not 4195GAT(1542) ; 4195GAT(1542)*
g3854 not 4251GAT(1566) ; 4251GAT(1566)*
g3855 not 4190GAT(1544) ; 4190GAT(1544)*
g3856 not 4248GAT(1567) ; 4248GAT(1567)*
g3857 not 4185GAT(1546) ; 4185GAT(1546)*
g3858 not 4245GAT(1568) ; 4245GAT(1568)*
g3859 not 4180GAT(1548) ; 4180GAT(1548)*
g3860 not 4242GAT(1570) ; 4242GAT(1570)*
g3861 not 4175GAT(1550) ; 4175GAT(1550)*
g3862 not 1296GAT(36) ; 1296GAT(36)*
g3863 not 4350GAT(1573) ; 4350GAT(1573)*
g3864 not 4348GAT(1574) ; 4348GAT(1574)*
g3865 not 4349GAT(1584) ; 4349GAT(1584)*
g3866 not 4344GAT(1585) ; 4344GAT(1585)*
g3867 not 4339GAT(1576) ; 4339GAT(1576)*
g3868 not 4340GAT(1577) ; 4340GAT(1577)*
g3869 not 4335GAT(1578) ; 4335GAT(1578)*
g3870 not 4332GAT(1579) ; 4332GAT(1579)*
g3871 not 4329GAT(1580) ; 4329GAT(1580)*
g3872 not 4327GAT(1581) ; 4327GAT(1581)*
g3873 not 4328GAT(1586) ; 4328GAT(1586)*
g3874 not 4323GAT(1587) ; 4323GAT(1587)*
g3875 not 4318GAT(1583) ; 4318GAT(1583)*
g3876 not 4319GAT(1588) ; 4319GAT(1588)*
g3877 not 4314GAT(1589) ; 4314GAT(1589)*
g3878 not 4310GAT(1590) ; 4310GAT(1590)*
g3879 not 4306GAT(1591) ; 4306GAT(1591)*
g3880 not 4341GAT(1575) ; 4341GAT(1575)*
g3881 not 1152GAT(84) ; 1152GAT(84)*
g3882 not 4302GAT(1592) ; 4302GAT(1592)*
g3883 not 4298GAT(1593) ; 4298GAT(1593)*
g3884 not 4294GAT(1594) ; 4294GAT(1594)*
g3885 not 4320GAT(1582) ; 4320GAT(1582)*
g3886 not 909GAT(165) ; 909GAT(165)*
g3887 not 4401GAT(1595) ; 4401GAT(1595)*
g3888 not 4398GAT(1596) ; 4398GAT(1596)*
g3889 not 4395GAT(1597) ; 4395GAT(1597)*
g3890 not 4393GAT(1598) ; 4393GAT(1598)*
g3891 not 4394GAT(1609) ; 4394GAT(1609)*
g3892 not 4389GAT(1611) ; 4389GAT(1611)*
g3893 not 4384GAT(1600) ; 4384GAT(1600)*
g3894 not 4385GAT(1601) ; 4385GAT(1601)*
g3895 not 4380GAT(1602) ; 4380GAT(1602)*
g3896 not 4377GAT(1603) ; 4377GAT(1603)*
g3897 not 4374GAT(1604) ; 4374GAT(1604)*
g3898 not 4372GAT(1605) ; 4372GAT(1605)*
g3899 not 4373GAT(1615) ; 4373GAT(1615)*
g3900 not 4368GAT(1616) ; 4368GAT(1616)*
g3901 not 4363GAT(1607) ; 4363GAT(1607)*
g3902 not 4364GAT(1617) ; 4364GAT(1617)*
g3903 not 4361GAT(1608) ; 4361GAT(1608)*
g3904 not 4362GAT(1618) ; 4362GAT(1618)*
g3905 not 4359GAT(1610) ; 4359GAT(1610)*
g3906 not 4360GAT(1619) ; 4360GAT(1619)*
g3907 not 4357GAT(1612) ; 4357GAT(1612)*
g3908 not 4358GAT(1620) ; 4358GAT(1620)*
g3909 not 4386GAT(1599) ; 4386GAT(1599)*
g3910 not 1104GAT(100) ; 1104GAT(100)*
g3911 not 4355GAT(1613) ; 4355GAT(1613)*
g3912 not 4356GAT(1621) ; 4356GAT(1621)*
g3913 not 4353GAT(1614) ; 4353GAT(1614)*
g3914 not 4354GAT(1622) ; 4354GAT(1622)*
g3915 not 4365GAT(1606) ; 4365GAT(1606)*
g3916 not 861GAT(181) ; 861GAT(181)*
g3917 not 4460GAT(1623) ; 4460GAT(1623)*
g3918 not 4461GAT(1624) ; 4461GAT(1624)*
g3919 not 4456GAT(1625) ; 4456GAT(1625)*
g3920 not 4453GAT(1626) ; 4453GAT(1626)*
g3921 not 4450GAT(1627) ; 4450GAT(1627)*
g3922 not 4448GAT(1628) ; 4448GAT(1628)*
g3923 not 4449GAT(1639) ; 4449GAT(1639)*
g3924 not 4444GAT(1641) ; 4444GAT(1641)*
g3925 not 4439GAT(1630) ; 4439GAT(1630)*
g3926 not 4440GAT(1631) ; 4440GAT(1631)*
g3927 not 4435GAT(1632) ; 4435GAT(1632)*
g3928 not 4432GAT(1633) ; 4432GAT(1633)*
g3929 not 4429GAT(1634) ; 4429GAT(1634)*
g3930 not 4427GAT(1635) ; 4427GAT(1635)*
g3931 not 4428GAT(1644) ; 4428GAT(1644)*
g3932 not 4423GAT(1645) ; 4423GAT(1645)*
g3933 not 4441GAT(1629) ; 4441GAT(1629)*
g3934 not 1056GAT(116) ; 1056GAT(116)*
g3935 not 4420GAT(1636) ; 4420GAT(1636)*
g3936 not 813GAT(197) ; 813GAT(197)*
g3937 not 4417GAT(1637) ; 4417GAT(1637)*
g3938 not 765GAT(213) ; 765GAT(213)*
g3939 not 4414GAT(1638) ; 4414GAT(1638)*
g3940 not 717GAT(229) ; 717GAT(229)*
g3941 not 4411GAT(1640) ; 4411GAT(1640)*
g3942 not 669GAT(245) ; 669GAT(245)*
g3943 not 4408GAT(1642) ; 4408GAT(1642)*
g3944 not 621GAT(261) ; 621GAT(261)*
g3945 not 4405GAT(1643) ; 4405GAT(1643)*
g3946 not 573GAT(277) ; 573GAT(277)*
g3947 not 4519GAT(1647) ; 4519GAT(1647)*
g3948 not 4520GAT(1648) ; 4520GAT(1648)*
g3949 not 4515GAT(1649) ; 4515GAT(1649)*
g3950 not 4512GAT(1650) ; 4512GAT(1650)*
g3951 not 4509GAT(1651) ; 4509GAT(1651)*
g3952 not 4507GAT(1652) ; 4507GAT(1652)*
g3953 not 4508GAT(1660) ; 4508GAT(1660)*
g3954 not 4503GAT(1661) ; 4503GAT(1661)*
g3955 not 4498GAT(1654) ; 4498GAT(1654)*
g3956 not 4499GAT(1655) ; 4499GAT(1655)*
g3957 not 4494GAT(1656) ; 4494GAT(1656)*
g3958 not 4491GAT(1657) ; 4491GAT(1657)*
g3959 not 4488GAT(1658) ; 4488GAT(1658)*
g3960 not 4486GAT(1659) ; 4486GAT(1659)*
g3961 not 4487GAT(1662) ; 4487GAT(1662)*
g3962 not 4482GAT(1663) ; 4482GAT(1663)*
g3963 not 4521GAT(1646) ; 4521GAT(1646)*
g3964 not 1251GAT(51) ; 1251GAT(51)*
g3965 not 4478GAT(1664) ; 4478GAT(1664)*
g3966 not 4474GAT(1665) ; 4474GAT(1665)*
g3967 not 4470GAT(1666) ; 4470GAT(1666)*
g3968 not 4466GAT(1667) ; 4466GAT(1667)*
g3969 not 4462GAT(1668) ; 4462GAT(1668)*
g3970 not 4500GAT(1653) ; 4500GAT(1653)*
g3971 not 1008GAT(132) ; 1008GAT(132)*
g3972 not 4587GAT(1682) ; 4587GAT(1682)*
g3973 not 4582GAT(1670) ; 4582GAT(1670)*
g3974 not 4583GAT(1671) ; 4583GAT(1671)*
g3975 not 4578GAT(1672) ; 4578GAT(1672)*
g3976 not 4575GAT(1673) ; 4575GAT(1673)*
g3977 not 4572GAT(1674) ; 4572GAT(1674)*
g3978 not 4570GAT(1675) ; 4570GAT(1675)*
g3979 not 4571GAT(1687) ; 4571GAT(1687)*
g3980 not 4566GAT(1689) ; 4566GAT(1689)*
g3981 not 4561GAT(1677) ; 4561GAT(1677)*
g3982 not 4562GAT(1678) ; 4562GAT(1678)*
g3983 not 4557GAT(1679) ; 4557GAT(1679)*
g3984 not 4554GAT(1680) ; 4554GAT(1680)*
g3985 not 4551GAT(1690) ; 4551GAT(1690)*
g3986 not 4549GAT(1681) ; 4549GAT(1681)*
g3987 not 4550GAT(1691) ; 4550GAT(1691)*
g3988 not 4544GAT(1683) ; 4544GAT(1683)*
g3989 not 4545GAT(1693) ; 4545GAT(1693)*
g3990 not 4584GAT(1669) ; 4584GAT(1669)*
g3991 not 1203GAT(67) ; 1203GAT(67)*
g3992 not 4539GAT(1684) ; 4539GAT(1684)*
g3993 not 4540GAT(1695) ; 4540GAT(1695)*
g3994 not 4534GAT(1685) ; 4534GAT(1685)*
g3995 not 4535GAT(1697) ; 4535GAT(1697)*
g3996 not 4529GAT(1686) ; 4529GAT(1686)*
g3997 not 4530GAT(1699) ; 4530GAT(1699)*
g3998 not 4524GAT(1688) ; 4524GAT(1688)*
g3999 not 4525GAT(1701) ; 4525GAT(1701)*
g4000 not 4563GAT(1676) ; 4563GAT(1676)*
g4001 not 960GAT(148) ; 960GAT(148)*
g4002 not 1299GAT(35) ; 1299GAT(35)*
g4003 not 4643GAT(1702) ; 4643GAT(1702)*
g4004 not 4641GAT(1703) ; 4641GAT(1703)*
g4005 not 4642GAT(1716) ; 4642GAT(1716)*
g4006 not 4637GAT(1718) ; 4637GAT(1718)*
g4007 not 4632GAT(1705) ; 4632GAT(1705)*
g4008 not 4633GAT(1706) ; 4633GAT(1706)*
g4009 not 4628GAT(1707) ; 4628GAT(1707)*
g4010 not 4625GAT(1708) ; 4625GAT(1708)*
g4011 not 4622GAT(1709) ; 4622GAT(1709)*
g4012 not 4620GAT(1710) ; 4620GAT(1710)*
g4013 not 4621GAT(1723) ; 4621GAT(1723)*
g4014 not 4616GAT(1724) ; 4616GAT(1724)*
g4015 not 4611GAT(1712) ; 4611GAT(1712)*
g4016 not 4612GAT(1713) ; 4612GAT(1713)*
g4017 not 4607GAT(1714) ; 4607GAT(1714)*
g4018 not 4634GAT(1704) ; 4634GAT(1704)*
g4019 not 1155GAT(83) ; 1155GAT(83)*
g4020 not 4613GAT(1711) ; 4613GAT(1711)*
g4021 not 912GAT(164) ; 912GAT(164)*
g4022 not 4604GAT(1715) ; 4604GAT(1715)*
g4023 not 4546GAT(1692) ; 4546GAT(1692)*
g4024 not 4601GAT(1717) ; 4601GAT(1717)*
g4025 not 4541GAT(1694) ; 4541GAT(1694)*
g4026 not 4598GAT(1719) ; 4598GAT(1719)*
g4027 not 4536GAT(1696) ; 4536GAT(1696)*
g4028 not 4595GAT(1720) ; 4595GAT(1720)*
g4029 not 4531GAT(1698) ; 4531GAT(1698)*
g4030 not 4592GAT(1721) ; 4592GAT(1721)*
g4031 not 4526GAT(1700) ; 4526GAT(1700)*
g4032 not 4704GAT(1725) ; 4704GAT(1725)*
g4033 not 4701GAT(1726) ; 4701GAT(1726)*
g4034 not 4698GAT(1727) ; 4698GAT(1727)*
g4035 not 4696GAT(1728) ; 4696GAT(1728)*
g4036 not 4697GAT(1738) ; 4697GAT(1738)*
g4037 not 4692GAT(1739) ; 4692GAT(1739)*
g4038 not 4687GAT(1730) ; 4687GAT(1730)*
g4039 not 4688GAT(1731) ; 4688GAT(1731)*
g4040 not 4683GAT(1732) ; 4683GAT(1732)*
g4041 not 4680GAT(1733) ; 4680GAT(1733)*
g4042 not 4677GAT(1734) ; 4677GAT(1734)*
g4043 not 4675GAT(1735) ; 4675GAT(1735)*
g4044 not 4676GAT(1740) ; 4676GAT(1740)*
g4045 not 4671GAT(1741) ; 4671GAT(1741)*
g4046 not 4666GAT(1737) ; 4666GAT(1737)*
g4047 not 4667GAT(1742) ; 4667GAT(1742)*
g4048 not 4662GAT(1743) ; 4662GAT(1743)*
g4049 not 4658GAT(1744) ; 4658GAT(1744)*
g4050 not 4654GAT(1745) ; 4654GAT(1745)*
g4051 not 4650GAT(1746) ; 4650GAT(1746)*
g4052 not 4689GAT(1729) ; 4689GAT(1729)*
g4053 not 1107GAT(99) ; 1107GAT(99)*
g4054 not 4646GAT(1747) ; 4646GAT(1747)*
g4055 not 4668GAT(1736) ; 4668GAT(1736)*
g4056 not 864GAT(180) ; 864GAT(180)*
g4057 not 4758GAT(1748) ; 4758GAT(1748)*
g4058 not 4759GAT(1749) ; 4759GAT(1749)*
g4059 not 4754GAT(1750) ; 4754GAT(1750)*
g4060 not 4751GAT(1751) ; 4751GAT(1751)*
g4061 not 4748GAT(1752) ; 4748GAT(1752)*
g4062 not 4746GAT(1753) ; 4746GAT(1753)*
g4063 not 4747GAT(1765) ; 4747GAT(1765)*
g4064 not 4742GAT(1767) ; 4742GAT(1767)*
g4065 not 4737GAT(1755) ; 4737GAT(1755)*
g4066 not 4738GAT(1756) ; 4738GAT(1756)*
g4067 not 4733GAT(1757) ; 4733GAT(1757)*
g4068 not 4730GAT(1758) ; 4730GAT(1758)*
g4069 not 4727GAT(1759) ; 4727GAT(1759)*
g4070 not 4725GAT(1760) ; 4725GAT(1760)*
g4071 not 4726GAT(1769) ; 4726GAT(1769)*
g4072 not 4721GAT(1770) ; 4721GAT(1770)*
g4073 not 4716GAT(1762) ; 4716GAT(1762)*
g4074 not 4717GAT(1771) ; 4717GAT(1771)*
g4075 not 4714GAT(1763) ; 4714GAT(1763)*
g4076 not 4715GAT(1772) ; 4715GAT(1772)*
g4077 not 4712GAT(1764) ; 4712GAT(1764)*
g4078 not 4713GAT(1773) ; 4713GAT(1773)*
g4079 not 4710GAT(1766) ; 4710GAT(1766)*
g4080 not 4711GAT(1774) ; 4711GAT(1774)*
g4081 not 4708GAT(1768) ; 4708GAT(1768)*
g4082 not 4709GAT(1775) ; 4709GAT(1775)*
g4083 not 4739GAT(1754) ; 4739GAT(1754)*
g4084 not 1059GAT(115) ; 1059GAT(115)*
g4085 not 4718GAT(1761) ; 4718GAT(1761)*
g4086 not 816GAT(196) ; 816GAT(196)*
g4087 not 4812GAT(1777) ; 4812GAT(1777)*
g4088 not 4813GAT(1778) ; 4813GAT(1778)*
g4089 not 4808GAT(1779) ; 4808GAT(1779)*
g4090 not 4805GAT(1780) ; 4805GAT(1780)*
g4091 not 4802GAT(1781) ; 4802GAT(1781)*
g4092 not 4800GAT(1782) ; 4800GAT(1782)*
g4093 not 4801GAT(1794) ; 4801GAT(1794)*
g4094 not 4796GAT(1796) ; 4796GAT(1796)*
g4095 not 4791GAT(1784) ; 4791GAT(1784)*
g4096 not 4792GAT(1785) ; 4792GAT(1785)*
g4097 not 4787GAT(1786) ; 4787GAT(1786)*
g4098 not 4784GAT(1787) ; 4784GAT(1787)*
g4099 not 4781GAT(1788) ; 4781GAT(1788)*
g4100 not 4779GAT(1789) ; 4779GAT(1789)*
g4101 not 4780GAT(1797) ; 4780GAT(1797)*
g4102 not 4775GAT(1798) ; 4775GAT(1798)*
g4103 not 4814GAT(1776) ; 4814GAT(1776)*
g4104 not 1254GAT(50) ; 1254GAT(50)*
g4105 not 4793GAT(1783) ; 4793GAT(1783)*
g4106 not 1011GAT(131) ; 1011GAT(131)*
g4107 not 4772GAT(1790) ; 4772GAT(1790)*
g4108 not 768GAT(212) ; 768GAT(212)*
g4109 not 4769GAT(1791) ; 4769GAT(1791)*
g4110 not 720GAT(228) ; 720GAT(228)*
g4111 not 4766GAT(1792) ; 4766GAT(1792)*
g4112 not 672GAT(244) ; 672GAT(244)*
g4113 not 4763GAT(1793) ; 4763GAT(1793)*
g4114 not 624GAT(260) ; 624GAT(260)*
g4115 not 4760GAT(1795) ; 4760GAT(1795)*
g4116 not 576GAT(276) ; 576GAT(276)*
g4117 not 4875GAT(1813) ; 4875GAT(1813)*
g4118 not 4870GAT(1800) ; 4870GAT(1800)*
g4119 not 4871GAT(1801) ; 4871GAT(1801)*
g4120 not 4866GAT(1802) ; 4866GAT(1802)*
g4121 not 4863GAT(1803) ; 4863GAT(1803)*
g4122 not 4860GAT(1804) ; 4860GAT(1804)*
g4123 not 4858GAT(1805) ; 4858GAT(1805)*
g4124 not 4859GAT(1814) ; 4859GAT(1814)*
g4125 not 4854GAT(1815) ; 4854GAT(1815)*
g4126 not 4849GAT(1807) ; 4849GAT(1807)*
g4127 not 4850GAT(1808) ; 4850GAT(1808)*
g4128 not 4845GAT(1809) ; 4845GAT(1809)*
g4129 not 4842GAT(1810) ; 4842GAT(1810)*
g4130 not 4839GAT(1811) ; 4839GAT(1811)*
g4131 not 4837GAT(1812) ; 4837GAT(1812)*
g4132 not 4838GAT(1816) ; 4838GAT(1816)*
g4133 not 4833GAT(1817) ; 4833GAT(1817)*
g4134 not 4829GAT(1818) ; 4829GAT(1818)*
g4135 not 4872GAT(1799) ; 4872GAT(1799)*
g4136 not 1206GAT(66) ; 1206GAT(66)*
g4137 not 4825GAT(1819) ; 4825GAT(1819)*
g4138 not 4821GAT(1820) ; 4821GAT(1820)*
g4139 not 4817GAT(1821) ; 4817GAT(1821)*
g4140 not 4851GAT(1806) ; 4851GAT(1806)*
g4141 not 963GAT(147) ; 963GAT(147)*
g4142 not 1302GAT(34) ; 1302GAT(34)*
g4143 not 4943GAT(1822) ; 4943GAT(1822)*
g4144 not 4941GAT(1823) ; 4941GAT(1823)*
g4145 not 4942GAT(1837) ; 4942GAT(1837)*
g4146 not 4937GAT(1839) ; 4937GAT(1839)*
g4147 not 4932GAT(1825) ; 4932GAT(1825)*
g4148 not 4933GAT(1826) ; 4933GAT(1826)*
g4149 not 4928GAT(1827) ; 4928GAT(1827)*
g4150 not 4925GAT(1828) ; 4925GAT(1828)*
g4151 not 4922GAT(1829) ; 4922GAT(1829)*
g4152 not 4920GAT(1830) ; 4920GAT(1830)*
g4153 not 4921GAT(1843) ; 4921GAT(1843)*
g4154 not 4916GAT(1844) ; 4916GAT(1844)*
g4155 not 4911GAT(1832) ; 4911GAT(1832)*
g4156 not 4912GAT(1833) ; 4912GAT(1833)*
g4157 not 4907GAT(1834) ; 4907GAT(1834)*
g4158 not 4904GAT(1835) ; 4904GAT(1835)*
g4159 not 4901GAT(1845) ; 4901GAT(1845)*
g4160 not 4899GAT(1836) ; 4899GAT(1836)*
g4161 not 4900GAT(1846) ; 4900GAT(1846)*
g4162 not 4894GAT(1838) ; 4894GAT(1838)*
g4163 not 4895GAT(1848) ; 4895GAT(1848)*
g4164 not 4889GAT(1840) ; 4889GAT(1840)*
g4165 not 4890GAT(1850) ; 4890GAT(1850)*
g4166 not 4934GAT(1824) ; 4934GAT(1824)*
g4167 not 1158GAT(82) ; 1158GAT(82)*
g4168 not 4884GAT(1841) ; 4884GAT(1841)*
g4169 not 4885GAT(1852) ; 4885GAT(1852)*
g4170 not 4879GAT(1842) ; 4879GAT(1842)*
g4171 not 4880GAT(1854) ; 4880GAT(1854)*
g4172 not 4913GAT(1831) ; 4913GAT(1831)*
g4173 not 915GAT(163) ; 915GAT(163)*
g4174 not 5001GAT(1855) ; 5001GAT(1855)*
g4175 not 4998GAT(1856) ; 4998GAT(1856)*
g4176 not 4995GAT(1857) ; 4995GAT(1857)*
g4177 not 4993GAT(1858) ; 4993GAT(1858)*
g4178 not 4994GAT(1872) ; 4994GAT(1872)*
g4179 not 4989GAT(1874) ; 4989GAT(1874)*
g4180 not 4984GAT(1860) ; 4984GAT(1860)*
g4181 not 4985GAT(1861) ; 4985GAT(1861)*
g4182 not 4980GAT(1862) ; 4980GAT(1862)*
g4183 not 4977GAT(1863) ; 4977GAT(1863)*
g4184 not 4974GAT(1864) ; 4974GAT(1864)*
g4185 not 4972GAT(1865) ; 4972GAT(1865)*
g4186 not 4973GAT(1877) ; 4973GAT(1877)*
g4187 not 4968GAT(1878) ; 4968GAT(1878)*
g4188 not 4963GAT(1867) ; 4963GAT(1867)*
g4189 not 4964GAT(1868) ; 4964GAT(1868)*
g4190 not 4959GAT(1869) ; 4959GAT(1869)*
g4191 not 4986GAT(1859) ; 4986GAT(1859)*
g4192 not 1110GAT(98) ; 1110GAT(98)*
g4193 not 4965GAT(1866) ; 4965GAT(1866)*
g4194 not 867GAT(179) ; 867GAT(179)*
g4195 not 4956GAT(1870) ; 4956GAT(1870)*
g4196 not 4896GAT(1847) ; 4896GAT(1847)*
g4197 not 4953GAT(1871) ; 4953GAT(1871)*
g4198 not 4891GAT(1849) ; 4891GAT(1849)*
g4199 not 4950GAT(1873) ; 4950GAT(1873)*
g4200 not 4886GAT(1851) ; 4886GAT(1851)*
g4201 not 4947GAT(1875) ; 4947GAT(1875)*
g4202 not 4881GAT(1853) ; 4881GAT(1853)*
g4203 not 5063GAT(1879) ; 5063GAT(1879)*
g4204 not 5064GAT(1880) ; 5064GAT(1880)*
g4205 not 5059GAT(1881) ; 5059GAT(1881)*
g4206 not 5056GAT(1882) ; 5056GAT(1882)*
g4207 not 5053GAT(1883) ; 5053GAT(1883)*
g4208 not 5051GAT(1884) ; 5051GAT(1884)*
g4209 not 5052GAT(1894) ; 5052GAT(1894)*
g4210 not 5047GAT(1895) ; 5047GAT(1895)*
g4211 not 5042GAT(1886) ; 5042GAT(1886)*
g4212 not 5043GAT(1887) ; 5043GAT(1887)*
g4213 not 5038GAT(1888) ; 5038GAT(1888)*
g4214 not 5035GAT(1889) ; 5035GAT(1889)*
g4215 not 5032GAT(1890) ; 5032GAT(1890)*
g4216 not 5030GAT(1891) ; 5030GAT(1891)*
g4217 not 5031GAT(1896) ; 5031GAT(1896)*
g4218 not 5026GAT(1897) ; 5026GAT(1897)*
g4219 not 5021GAT(1893) ; 5021GAT(1893)*
g4220 not 5022GAT(1898) ; 5022GAT(1898)*
g4221 not 5017GAT(1899) ; 5017GAT(1899)*
g4222 not 5013GAT(1900) ; 5013GAT(1900)*
g4223 not 5009GAT(1901) ; 5009GAT(1901)*
g4224 not 5005GAT(1902) ; 5005GAT(1902)*
g4225 not 5044GAT(1885) ; 5044GAT(1885)*
g4226 not 1062GAT(114) ; 1062GAT(114)*
g4227 not 5023GAT(1892) ; 5023GAT(1892)*
g4228 not 819GAT(195) ; 819GAT(195)*
g4229 not 5113GAT(1904) ; 5113GAT(1904)*
g4230 not 5114GAT(1905) ; 5114GAT(1905)*
g4231 not 5109GAT(1906) ; 5109GAT(1906)*
g4232 not 5106GAT(1907) ; 5106GAT(1907)*
g4233 not 5103GAT(1908) ; 5103GAT(1908)*
g4234 not 5101GAT(1909) ; 5101GAT(1909)*
g4235 not 5102GAT(1922) ; 5102GAT(1922)*
g4236 not 5097GAT(1923) ; 5097GAT(1923)*
g4237 not 5092GAT(1911) ; 5092GAT(1911)*
g4238 not 5093GAT(1912) ; 5093GAT(1912)*
g4239 not 5088GAT(1913) ; 5088GAT(1913)*
g4240 not 5085GAT(1914) ; 5085GAT(1914)*
g4241 not 5082GAT(1915) ; 5082GAT(1915)*
g4242 not 5080GAT(1916) ; 5080GAT(1916)*
g4243 not 5081GAT(1924) ; 5081GAT(1924)*
g4244 not 5076GAT(1925) ; 5076GAT(1925)*
g4245 not 5071GAT(1918) ; 5071GAT(1918)*
g4246 not 5072GAT(1926) ; 5072GAT(1926)*
g4247 not 5115GAT(1903) ; 5115GAT(1903)*
g4248 not 1257GAT(49) ; 1257GAT(49)*
g4249 not 5069GAT(1919) ; 5069GAT(1919)*
g4250 not 5070GAT(1927) ; 5070GAT(1927)*
g4251 not 5067GAT(1920) ; 5067GAT(1920)*
g4252 not 5068GAT(1928) ; 5068GAT(1928)*
g4253 not 5065GAT(1921) ; 5065GAT(1921)*
g4254 not 5066GAT(1929) ; 5066GAT(1929)*
g4255 not 5094GAT(1910) ; 5094GAT(1910)*
g4256 not 1014GAT(130) ; 1014GAT(130)*
g4257 not 5073GAT(1917) ; 5073GAT(1917)*
g4258 not 771GAT(211) ; 771GAT(211)*
g4259 not 5172GAT(1945) ; 5172GAT(1945)*
g4260 not 5167GAT(1931) ; 5167GAT(1931)*
g4261 not 5168GAT(1932) ; 5168GAT(1932)*
g4262 not 5163GAT(1933) ; 5163GAT(1933)*
g4263 not 5160GAT(1934) ; 5160GAT(1934)*
g4264 not 5157GAT(1935) ; 5157GAT(1935)*
g4265 not 5155GAT(1936) ; 5155GAT(1936)*
g4266 not 5156GAT(1949) ; 5156GAT(1949)*
g4267 not 5151GAT(1950) ; 5151GAT(1950)*
g4268 not 5146GAT(1938) ; 5146GAT(1938)*
g4269 not 5147GAT(1939) ; 5147GAT(1939)*
g4270 not 5142GAT(1940) ; 5142GAT(1940)*
g4271 not 5139GAT(1941) ; 5139GAT(1941)*
g4272 not 5136GAT(1942) ; 5136GAT(1942)*
g4273 not 5134GAT(1943) ; 5134GAT(1943)*
g4274 not 5135GAT(1951) ; 5135GAT(1951)*
g4275 not 5130GAT(1952) ; 5130GAT(1952)*
g4276 not 5169GAT(1930) ; 5169GAT(1930)*
g4277 not 1209GAT(65) ; 1209GAT(65)*
g4278 not 5148GAT(1937) ; 5148GAT(1937)*
g4279 not 966GAT(146) ; 966GAT(146)*
g4280 not 5127GAT(1944) ; 5127GAT(1944)*
g4281 not 723GAT(227) ; 723GAT(227)*
g4282 not 5124GAT(1946) ; 5124GAT(1946)*
g4283 not 675GAT(243) ; 675GAT(243)*
g4284 not 5121GAT(1947) ; 5121GAT(1947)*
g4285 not 627GAT(259) ; 627GAT(259)*
g4286 not 5118GAT(1948) ; 5118GAT(1948)*
g4287 not 579GAT(275) ; 579GAT(275)*
g4288 not 1305GAT(33) ; 1305GAT(33)*
g4289 not 5236GAT(1953) ; 5236GAT(1953)*
g4290 not 5234GAT(1954) ; 5234GAT(1954)*
g4291 not 5235GAT(1969) ; 5235GAT(1969)*
g4292 not 5230GAT(1970) ; 5230GAT(1970)*
g4293 not 5225GAT(1956) ; 5225GAT(1956)*
g4294 not 5226GAT(1957) ; 5226GAT(1957)*
g4295 not 5221GAT(1958) ; 5221GAT(1958)*
g4296 not 5218GAT(1959) ; 5218GAT(1959)*
g4297 not 5215GAT(1960) ; 5215GAT(1960)*
g4298 not 5213GAT(1961) ; 5213GAT(1961)*
g4299 not 5214GAT(1971) ; 5214GAT(1971)*
g4300 not 5209GAT(1972) ; 5209GAT(1972)*
g4301 not 5204GAT(1963) ; 5204GAT(1963)*
g4302 not 5205GAT(1964) ; 5205GAT(1964)*
g4303 not 5200GAT(1965) ; 5200GAT(1965)*
g4304 not 5197GAT(1966) ; 5197GAT(1966)*
g4305 not 5194GAT(1967) ; 5194GAT(1967)*
g4306 not 5192GAT(1968) ; 5192GAT(1968)*
g4307 not 5193GAT(1973) ; 5193GAT(1973)*
g4308 not 5188GAT(1974) ; 5188GAT(1974)*
g4309 not 5184GAT(1975) ; 5184GAT(1975)*
g4310 not 5180GAT(1976) ; 5180GAT(1976)*
g4311 not 5227GAT(1955) ; 5227GAT(1955)*
g4312 not 1161GAT(81) ; 1161GAT(81)*
g4313 not 5176GAT(1977) ; 5176GAT(1977)*
g4314 not 5206GAT(1962) ; 5206GAT(1962)*
g4315 not 918GAT(162) ; 918GAT(162)*
g4316 not 5304GAT(1978) ; 5304GAT(1978)*
g4317 not 5301GAT(1979) ; 5301GAT(1979)*
g4318 not 5298GAT(1980) ; 5298GAT(1980)*
g4319 not 5296GAT(1981) ; 5296GAT(1981)*
g4320 not 5297GAT(1996) ; 5297GAT(1996)*
g4321 not 5292GAT(1998) ; 5292GAT(1998)*
g4322 not 5287GAT(1983) ; 5287GAT(1983)*
g4323 not 5288GAT(1984) ; 5288GAT(1984)*
g4324 not 5283GAT(1985) ; 5283GAT(1985)*
g4325 not 5280GAT(1986) ; 5280GAT(1986)*
g4326 not 5277GAT(1987) ; 5277GAT(1987)*
g4327 not 5275GAT(1988) ; 5275GAT(1988)*
g4328 not 5276GAT(2000) ; 5276GAT(2000)*
g4329 not 5271GAT(2001) ; 5271GAT(2001)*
g4330 not 5266GAT(1990) ; 5266GAT(1990)*
g4331 not 5267GAT(1991) ; 5267GAT(1991)*
g4332 not 5262GAT(1992) ; 5262GAT(1992)*
g4333 not 5259GAT(1993) ; 5259GAT(1993)*
g4334 not 5256GAT(2002) ; 5256GAT(2002)*
g4335 not 5254GAT(1994) ; 5254GAT(1994)*
g4336 not 5255GAT(2003) ; 5255GAT(2003)*
g4337 not 5249GAT(1995) ; 5249GAT(1995)*
g4338 not 5250GAT(2005) ; 5250GAT(2005)*
g4339 not 5244GAT(1997) ; 5244GAT(1997)*
g4340 not 5245GAT(2007) ; 5245GAT(2007)*
g4341 not 5239GAT(1999) ; 5239GAT(1999)*
g4342 not 5240GAT(2009) ; 5240GAT(2009)*
g4343 not 5289GAT(1982) ; 5289GAT(1982)*
g4344 not 1113GAT(97) ; 1113GAT(97)*
g4345 not 5268GAT(1989) ; 5268GAT(1989)*
g4346 not 870GAT(178) ; 870GAT(178)*
g4347 not 5364GAT(2010) ; 5364GAT(2010)*
g4348 not 5365GAT(2011) ; 5365GAT(2011)*
g4349 not 5360GAT(2012) ; 5360GAT(2012)*
g4350 not 5357GAT(2013) ; 5357GAT(2013)*
g4351 not 5354GAT(2014) ; 5354GAT(2014)*
g4352 not 5352GAT(2015) ; 5352GAT(2015)*
g4353 not 5353GAT(2030) ; 5353GAT(2030)*
g4354 not 5348GAT(2032) ; 5348GAT(2032)*
g4355 not 5343GAT(2017) ; 5343GAT(2017)*
g4356 not 5344GAT(2018) ; 5344GAT(2018)*
g4357 not 5339GAT(2019) ; 5339GAT(2019)*
g4358 not 5336GAT(2020) ; 5336GAT(2020)*
g4359 not 5333GAT(2021) ; 5333GAT(2021)*
g4360 not 5331GAT(2022) ; 5331GAT(2022)*
g4361 not 5332GAT(2033) ; 5332GAT(2033)*
g4362 not 5327GAT(2034) ; 5327GAT(2034)*
g4363 not 5322GAT(2024) ; 5322GAT(2024)*
g4364 not 5323GAT(2025) ; 5323GAT(2025)*
g4365 not 5318GAT(2026) ; 5318GAT(2026)*
g4366 not 5345GAT(2016) ; 5345GAT(2016)*
g4367 not 1065GAT(113) ; 1065GAT(113)*
g4368 not 5324GAT(2023) ; 5324GAT(2023)*
g4369 not 822GAT(194) ; 822GAT(194)*
g4370 not 5315GAT(2027) ; 5315GAT(2027)*
g4371 not 5251GAT(2004) ; 5251GAT(2004)*
g4372 not 5312GAT(2028) ; 5312GAT(2028)*
g4373 not 5246GAT(2006) ; 5246GAT(2006)*
g4374 not 5309GAT(2029) ; 5309GAT(2029)*
g4375 not 5241GAT(2008) ; 5241GAT(2008)*
g4376 not 5420GAT(2036) ; 5420GAT(2036)*
g4377 not 5421GAT(2037) ; 5421GAT(2037)*
g4378 not 5416GAT(2038) ; 5416GAT(2038)*
g4379 not 5413GAT(2039) ; 5413GAT(2039)*
g4380 not 5410GAT(2040) ; 5410GAT(2040)*
g4381 not 5408GAT(2041) ; 5408GAT(2041)*
g4382 not 5409GAT(2051) ; 5409GAT(2051)*
g4383 not 5404GAT(2052) ; 5404GAT(2052)*
g4384 not 5399GAT(2043) ; 5399GAT(2043)*
g4385 not 5400GAT(2044) ; 5400GAT(2044)*
g4386 not 5395GAT(2045) ; 5395GAT(2045)*
g4387 not 5392GAT(2046) ; 5392GAT(2046)*
g4388 not 5389GAT(2047) ; 5389GAT(2047)*
g4389 not 5387GAT(2048) ; 5387GAT(2048)*
g4390 not 5388GAT(2053) ; 5388GAT(2053)*
g4391 not 5383GAT(2054) ; 5383GAT(2054)*
g4392 not 5378GAT(2050) ; 5378GAT(2050)*
g4393 not 5379GAT(2055) ; 5379GAT(2055)*
g4394 not 5374GAT(2056) ; 5374GAT(2056)*
g4395 not 5422GAT(2035) ; 5422GAT(2035)*
g4396 not 1260GAT(48) ; 1260GAT(48)*
g4397 not 5370GAT(2057) ; 5370GAT(2057)*
g4398 not 5366GAT(2058) ; 5366GAT(2058)*
g4399 not 5401GAT(2042) ; 5401GAT(2042)*
g4400 not 1017GAT(129) ; 1017GAT(129)*
g4401 not 5380GAT(2049) ; 5380GAT(2049)*
g4402 not 774GAT(210) ; 774GAT(210)*
g4403 not 5476GAT(2075) ; 5476GAT(2075)*
g4404 not 5471GAT(2060) ; 5471GAT(2060)*
g4405 not 5472GAT(2061) ; 5472GAT(2061)*
g4406 not 5467GAT(2062) ; 5467GAT(2062)*
g4407 not 5464GAT(2063) ; 5464GAT(2063)*
g4408 not 5461GAT(2064) ; 5461GAT(2064)*
g4409 not 5459GAT(2065) ; 5459GAT(2065)*
g4410 not 5460GAT(2078) ; 5460GAT(2078)*
g4411 not 5455GAT(2079) ; 5455GAT(2079)*
g4412 not 5450GAT(2067) ; 5450GAT(2067)*
g4413 not 5451GAT(2068) ; 5451GAT(2068)*
g4414 not 5446GAT(2069) ; 5446GAT(2069)*
g4415 not 5443GAT(2070) ; 5443GAT(2070)*
g4416 not 5440GAT(2071) ; 5440GAT(2071)*
g4417 not 5438GAT(2072) ; 5438GAT(2072)*
g4418 not 5439GAT(2080) ; 5439GAT(2080)*
g4419 not 5434GAT(2081) ; 5434GAT(2081)*
g4420 not 5429GAT(2074) ; 5429GAT(2074)*
g4421 not 5430GAT(2082) ; 5430GAT(2082)*
g4422 not 5427GAT(2076) ; 5427GAT(2076)*
g4423 not 5428GAT(2083) ; 5428GAT(2083)*
g4424 not 5473GAT(2059) ; 5473GAT(2059)*
g4425 not 1212GAT(64) ; 1212GAT(64)*
g4426 not 5425GAT(2077) ; 5425GAT(2077)*
g4427 not 5426GAT(2084) ; 5426GAT(2084)*
g4428 not 5452GAT(2066) ; 5452GAT(2066)*
g4429 not 969GAT(145) ; 969GAT(145)*
g4430 not 5431GAT(2073) ; 5431GAT(2073)*
g4431 not 726GAT(226) ; 726GAT(226)*
g4432 not 1308GAT(32) ; 1308GAT(32)*
g4433 not 5537GAT(2085) ; 5537GAT(2085)*
g4434 not 5535GAT(2086) ; 5535GAT(2086)*
g4435 not 5536GAT(2102) ; 5536GAT(2102)*
g4436 not 5531GAT(2104) ; 5531GAT(2104)*
g4437 not 5526GAT(2088) ; 5526GAT(2088)*
g4438 not 5527GAT(2089) ; 5527GAT(2089)*
g4439 not 5522GAT(2090) ; 5522GAT(2090)*
g4440 not 5519GAT(2091) ; 5519GAT(2091)*
g4441 not 5516GAT(2092) ; 5516GAT(2092)*
g4442 not 5514GAT(2093) ; 5514GAT(2093)*
g4443 not 5515GAT(2106) ; 5515GAT(2106)*
g4444 not 5510GAT(2107) ; 5510GAT(2107)*
g4445 not 5505GAT(2095) ; 5505GAT(2095)*
g4446 not 5506GAT(2096) ; 5506GAT(2096)*
g4447 not 5501GAT(2097) ; 5501GAT(2097)*
g4448 not 5498GAT(2098) ; 5498GAT(2098)*
g4449 not 5495GAT(2099) ; 5495GAT(2099)*
g4450 not 5493GAT(2100) ; 5493GAT(2100)*
g4451 not 5494GAT(2108) ; 5494GAT(2108)*
g4452 not 5489GAT(2109) ; 5489GAT(2109)*
g4453 not 5528GAT(2087) ; 5528GAT(2087)*
g4454 not 1164GAT(80) ; 1164GAT(80)*
g4455 not 5507GAT(2094) ; 5507GAT(2094)*
g4456 not 921GAT(161) ; 921GAT(161)*
g4457 not 5486GAT(2101) ; 5486GAT(2101)*
g4458 not 678GAT(242) ; 678GAT(242)*
g4459 not 5483GAT(2103) ; 5483GAT(2103)*
g4460 not 630GAT(258) ; 630GAT(258)*
g4461 not 5480GAT(2105) ; 5480GAT(2105)*
g4462 not 582GAT(274) ; 582GAT(274)*
g4463 not 5602GAT(2110) ; 5602GAT(2110)*
g4464 not 5599GAT(2111) ; 5599GAT(2111)*
g4465 not 5596GAT(2112) ; 5596GAT(2112)*
g4466 not 5594GAT(2113) ; 5594GAT(2113)*
g4467 not 5595GAT(2128) ; 5595GAT(2128)*
g4468 not 5590GAT(2129) ; 5590GAT(2129)*
g4469 not 5585GAT(2115) ; 5585GAT(2115)*
g4470 not 5586GAT(2116) ; 5586GAT(2116)*
g4471 not 5581GAT(2117) ; 5581GAT(2117)*
g4472 not 5578GAT(2118) ; 5578GAT(2118)*
g4473 not 5575GAT(2119) ; 5575GAT(2119)*
g4474 not 5573GAT(2120) ; 5573GAT(2120)*
g4475 not 5574GAT(2130) ; 5574GAT(2130)*
g4476 not 5569GAT(2131) ; 5569GAT(2131)*
g4477 not 5564GAT(2122) ; 5564GAT(2122)*
g4478 not 5565GAT(2123) ; 5565GAT(2123)*
g4479 not 5560GAT(2124) ; 5560GAT(2124)*
g4480 not 5557GAT(2125) ; 5557GAT(2125)*
g4481 not 5554GAT(2126) ; 5554GAT(2126)*
g4482 not 5552GAT(2127) ; 5552GAT(2127)*
g4483 not 5553GAT(2132) ; 5553GAT(2132)*
g4484 not 5548GAT(2133) ; 5548GAT(2133)*
g4485 not 5544GAT(2134) ; 5544GAT(2134)*
g4486 not 5540GAT(2135) ; 5540GAT(2135)*
g4487 not 5587GAT(2114) ; 5587GAT(2114)*
g4488 not 1116GAT(96) ; 1116GAT(96)*
g4489 not 5566GAT(2121) ; 5566GAT(2121)*
g4490 not 873GAT(177) ; 873GAT(177)*
g4491 not 5670GAT(2136) ; 5670GAT(2136)*
g4492 not 5671GAT(2137) ; 5671GAT(2137)*
g4493 not 5666GAT(2138) ; 5666GAT(2138)*
g4494 not 5663GAT(2139) ; 5663GAT(2139)*
g4495 not 5660GAT(2140) ; 5660GAT(2140)*
g4496 not 5658GAT(2141) ; 5658GAT(2141)*
g4497 not 5659GAT(2157) ; 5659GAT(2157)*
g4498 not 5654GAT(2158) ; 5654GAT(2158)*
g4499 not 5649GAT(2143) ; 5649GAT(2143)*
g4500 not 5650GAT(2144) ; 5650GAT(2144)*
g4501 not 5645GAT(2145) ; 5645GAT(2145)*
g4502 not 5642GAT(2146) ; 5642GAT(2146)*
g4503 not 5639GAT(2147) ; 5639GAT(2147)*
g4504 not 5637GAT(2148) ; 5637GAT(2148)*
g4505 not 5638GAT(2159) ; 5638GAT(2159)*
g4506 not 5633GAT(2160) ; 5633GAT(2160)*
g4507 not 5628GAT(2150) ; 5628GAT(2150)*
g4508 not 5629GAT(2151) ; 5629GAT(2151)*
g4509 not 5624GAT(2152) ; 5624GAT(2152)*
g4510 not 5621GAT(2153) ; 5621GAT(2153)*
g4511 not 5618GAT(2161) ; 5618GAT(2161)*
g4512 not 5616GAT(2154) ; 5616GAT(2154)*
g4513 not 5617GAT(2162) ; 5617GAT(2162)*
g4514 not 5611GAT(2155) ; 5611GAT(2155)*
g4515 not 5612GAT(2164) ; 5612GAT(2164)*
g4516 not 5606GAT(2156) ; 5606GAT(2156)*
g4517 not 5607GAT(2166) ; 5607GAT(2166)*
g4518 not 5651GAT(2142) ; 5651GAT(2142)*
g4519 not 1068GAT(112) ; 1068GAT(112)*
g4520 not 5630GAT(2149) ; 5630GAT(2149)*
g4521 not 825GAT(193) ; 825GAT(193)*
g4522 not 5725GAT(2168) ; 5725GAT(2168)*
g4523 not 5726GAT(2169) ; 5726GAT(2169)*
g4524 not 5721GAT(2170) ; 5721GAT(2170)*
g4525 not 5718GAT(2171) ; 5718GAT(2171)*
g4526 not 5715GAT(2172) ; 5715GAT(2172)*
g4527 not 5713GAT(2173) ; 5713GAT(2173)*
g4528 not 5714GAT(2188) ; 5714GAT(2188)*
g4529 not 5709GAT(2189) ; 5709GAT(2189)*
g4530 not 5704GAT(2175) ; 5704GAT(2175)*
g4531 not 5705GAT(2176) ; 5705GAT(2176)*
g4532 not 5700GAT(2177) ; 5700GAT(2177)*
g4533 not 5697GAT(2178) ; 5697GAT(2178)*
g4534 not 5694GAT(2179) ; 5694GAT(2179)*
g4535 not 5692GAT(2180) ; 5692GAT(2180)*
g4536 not 5693GAT(2190) ; 5693GAT(2190)*
g4537 not 5688GAT(2191) ; 5688GAT(2191)*
g4538 not 5683GAT(2182) ; 5683GAT(2182)*
g4539 not 5684GAT(2183) ; 5684GAT(2183)*
g4540 not 5679GAT(2184) ; 5679GAT(2184)*
g4541 not 5706GAT(2174) ; 5706GAT(2174)*
g4542 not 1020GAT(128) ; 1020GAT(128)*
g4543 not 5685GAT(2181) ; 5685GAT(2181)*
g4544 not 777GAT(209) ; 777GAT(209)*
g4545 not 5676GAT(2185) ; 5676GAT(2185)*
g4546 not 5613GAT(2163) ; 5613GAT(2163)*
g4547 not 5673GAT(2186) ; 5673GAT(2186)*
g4548 not 5608GAT(2165) ; 5608GAT(2165)*
g4549 not 5780GAT(2193) ; 5780GAT(2193)*
g4550 not 5781GAT(2194) ; 5781GAT(2194)*
g4551 not 5776GAT(2195) ; 5776GAT(2195)*
g4552 not 5773GAT(2196) ; 5773GAT(2196)*
g4553 not 5770GAT(2197) ; 5770GAT(2197)*
g4554 not 5768GAT(2198) ; 5768GAT(2198)*
g4555 not 5769GAT(2208) ; 5769GAT(2208)*
g4556 not 5764GAT(2209) ; 5764GAT(2209)*
g4557 not 5759GAT(2200) ; 5759GAT(2200)*
g4558 not 5760GAT(2201) ; 5760GAT(2201)*
g4559 not 5755GAT(2202) ; 5755GAT(2202)*
g4560 not 5752GAT(2203) ; 5752GAT(2203)*
g4561 not 5749GAT(2204) ; 5749GAT(2204)*
g4562 not 5747GAT(2205) ; 5747GAT(2205)*
g4563 not 5748GAT(2210) ; 5748GAT(2210)*
g4564 not 5743GAT(2211) ; 5743GAT(2211)*
g4565 not 5738GAT(2207) ; 5738GAT(2207)*
g4566 not 5739GAT(2212) ; 5739GAT(2212)*
g4567 not 5734GAT(2213) ; 5734GAT(2213)*
g4568 not 5730GAT(2214) ; 5730GAT(2214)*
g4569 not 5761GAT(2199) ; 5761GAT(2199)*
g4570 not 972GAT(144) ; 972GAT(144)*
g4571 not 5740GAT(2206) ; 5740GAT(2206)*
g4572 not 729GAT(225) ; 729GAT(225)*
g4573 not 5829GAT(2216) ; 5829GAT(2216)*
g4574 not 5830GAT(2217) ; 5830GAT(2217)*
g4575 not 5825GAT(2218) ; 5825GAT(2218)*
g4576 not 5822GAT(2219) ; 5822GAT(2219)*
g4577 not 5819GAT(2220) ; 5819GAT(2220)*
g4578 not 5817GAT(2221) ; 5817GAT(2221)*
g4579 not 5818GAT(2232) ; 5818GAT(2232)*
g4580 not 5813GAT(2233) ; 5813GAT(2233)*
g4581 not 5808GAT(2223) ; 5808GAT(2223)*
g4582 not 5809GAT(2224) ; 5809GAT(2224)*
g4583 not 5804GAT(2225) ; 5804GAT(2225)*
g4584 not 5801GAT(2226) ; 5801GAT(2226)*
g4585 not 5798GAT(2227) ; 5798GAT(2227)*
g4586 not 5796GAT(2228) ; 5796GAT(2228)*
g4587 not 5797GAT(2234) ; 5797GAT(2234)*
g4588 not 5792GAT(2235) ; 5792GAT(2235)*
g4589 not 5787GAT(2230) ; 5787GAT(2230)*
g4590 not 5788GAT(2236) ; 5788GAT(2236)*
g4591 not 5785GAT(2231) ; 5785GAT(2231)*
g4592 not 5786GAT(2237) ; 5786GAT(2237)*
g4593 not 5810GAT(2222) ; 5810GAT(2222)*
g4594 not 924GAT(160) ; 924GAT(160)*
g4595 not 5789GAT(2229) ; 5789GAT(2229)*
g4596 not 681GAT(241) ; 681GAT(241)*
g4597 not 5877GAT(2239) ; 5877GAT(2239)*
g4598 not 5878GAT(2240) ; 5878GAT(2240)*
g4599 not 5873GAT(2241) ; 5873GAT(2241)*
g4600 not 5870GAT(2242) ; 5870GAT(2242)*
g4601 not 5867GAT(2243) ; 5867GAT(2243)*
g4602 not 5865GAT(2244) ; 5865GAT(2244)*
g4603 not 5866GAT(2254) ; 5866GAT(2254)*
g4604 not 5861GAT(2255) ; 5861GAT(2255)*
g4605 not 5856GAT(2246) ; 5856GAT(2246)*
g4606 not 5857GAT(2247) ; 5857GAT(2247)*
g4607 not 5852GAT(2248) ; 5852GAT(2248)*
g4608 not 5849GAT(2249) ; 5849GAT(2249)*
g4609 not 5846GAT(2250) ; 5846GAT(2250)*
g4610 not 5844GAT(2251) ; 5844GAT(2251)*
g4611 not 5845GAT(2256) ; 5845GAT(2256)*
g4612 not 5840GAT(2257) ; 5840GAT(2257)*
g4613 not 5858GAT(2245) ; 5858GAT(2245)*
g4614 not 876GAT(176) ; 876GAT(176)*
g4615 not 5837GAT(2252) ; 5837GAT(2252)*
g4616 not 633GAT(257) ; 633GAT(257)*
g4617 not 5834GAT(2253) ; 5834GAT(2253)*
g4618 not 585GAT(273) ; 585GAT(273)*
g4619 not 5923GAT(2259) ; 5923GAT(2259)*
g4620 not 5924GAT(2260) ; 5924GAT(2260)*
g4621 not 5919GAT(2261) ; 5919GAT(2261)*
g4622 not 5916GAT(2262) ; 5916GAT(2262)*
g4623 not 5913GAT(2263) ; 5913GAT(2263)*
g4624 not 5911GAT(2264) ; 5911GAT(2264)*
g4625 not 5912GAT(2272) ; 5912GAT(2272)*
g4626 not 5907GAT(2273) ; 5907GAT(2273)*
g4627 not 5902GAT(2266) ; 5902GAT(2266)*
g4628 not 5903GAT(2267) ; 5903GAT(2267)*
g4629 not 5898GAT(2268) ; 5898GAT(2268)*
g4630 not 5895GAT(2269) ; 5895GAT(2269)*
g4631 not 5892GAT(2270) ; 5892GAT(2270)*
g4632 not 5890GAT(2271) ; 5890GAT(2271)*
g4633 not 5891GAT(2274) ; 5891GAT(2274)*
g4634 not 5886GAT(2275) ; 5886GAT(2275)*
g4635 not 5882GAT(2276) ; 5882GAT(2276)*
g4636 not 5904GAT(2265) ; 5904GAT(2265)*
g4637 not 828GAT(192) ; 828GAT(192)*
g4638 not 5966GAT(2278) ; 5966GAT(2278)*
g4639 not 5967GAT(2279) ; 5967GAT(2279)*
g4640 not 5962GAT(2280) ; 5962GAT(2280)*
g4641 not 5959GAT(2281) ; 5959GAT(2281)*
g4642 not 5956GAT(2282) ; 5956GAT(2282)*
g4643 not 5954GAT(2283) ; 5954GAT(2283)*
g4644 not 5955GAT(2291) ; 5955GAT(2291)*
g4645 not 5950GAT(2292) ; 5950GAT(2292)*
g4646 not 5945GAT(2285) ; 5945GAT(2285)*
g4647 not 5946GAT(2286) ; 5946GAT(2286)*
g4648 not 5941GAT(2287) ; 5941GAT(2287)*
g4649 not 5938GAT(2288) ; 5938GAT(2288)*
g4650 not 5935GAT(2293) ; 5935GAT(2293)*
g4651 not 5933GAT(2289) ; 5933GAT(2289)*
g4652 not 5934GAT(2294) ; 5934GAT(2294)*
g4653 not 5928GAT(2290) ; 5928GAT(2290)*
g4654 not 5929GAT(2296) ; 5929GAT(2296)*
g4655 not 5947GAT(2284) ; 5947GAT(2284)*
g4656 not 780GAT(208) ; 780GAT(208)*
g4657 not 6000GAT(2298) ; 6000GAT(2298)*
g4658 not 6001GAT(2299) ; 6001GAT(2299)*
g4659 not 5996GAT(2300) ; 5996GAT(2300)*
g4660 not 5993GAT(2301) ; 5993GAT(2301)*
g4661 not 5990GAT(2302) ; 5990GAT(2302)*
g4662 not 5988GAT(2303) ; 5988GAT(2303)*
g4663 not 5989GAT(2310) ; 5989GAT(2310)*
g4664 not 5984GAT(2311) ; 5984GAT(2311)*
g4665 not 5979GAT(2305) ; 5979GAT(2305)*
g4666 not 5980GAT(2306) ; 5980GAT(2306)*
g4667 not 5975GAT(2307) ; 5975GAT(2307)*
g4668 not 5981GAT(2304) ; 5981GAT(2304)*
g4669 not 732GAT(224) ; 732GAT(224)*
g4670 not 5972GAT(2308) ; 5972GAT(2308)*
g4671 not 5930GAT(2295) ; 5930GAT(2295)*
g4672 not 6030GAT(2313) ; 6030GAT(2313)*
g4673 not 6031GAT(2314) ; 6031GAT(2314)*
g4674 not 6026GAT(2315) ; 6026GAT(2315)*
g4675 not 6023GAT(2316) ; 6023GAT(2316)*
g4676 not 6020GAT(2317) ; 6020GAT(2317)*
g4677 not 6018GAT(2318) ; 6018GAT(2318)*
g4678 not 6019GAT(2321) ; 6019GAT(2321)*
g4679 not 6014GAT(2322) ; 6014GAT(2322)*
g4680 not 6009GAT(2320) ; 6009GAT(2320)*
g4681 not 6010GAT(2323) ; 6010GAT(2323)*
g4682 not 6005GAT(2324) ; 6005GAT(2324)*
g4683 not 6011GAT(2319) ; 6011GAT(2319)*
g4684 not 684GAT(240) ; 684GAT(240)*
g4685 not 6056GAT(2326) ; 6056GAT(2326)*
g4686 not 6057GAT(2327) ; 6057GAT(2327)*
g4687 not 6052GAT(2328) ; 6052GAT(2328)*
g4688 not 6049GAT(2329) ; 6049GAT(2329)*
g4689 not 6046GAT(2330) ; 6046GAT(2330)*
g4690 not 6044GAT(2331) ; 6044GAT(2331)*
g4691 not 6045GAT(2334) ; 6045GAT(2334)*
g4692 not 6040GAT(2335) ; 6040GAT(2335)*
g4693 not 6035GAT(2333) ; 6035GAT(2333)*
g4694 not 6036GAT(2336) ; 6036GAT(2336)*
g4695 not 6037GAT(2332) ; 6037GAT(2332)*
g4696 not 636GAT(256) ; 636GAT(256)*
g4697 not 6080GAT(2338) ; 6080GAT(2338)*
g4698 not 6081GAT(2339) ; 6081GAT(2339)*
g4699 not 6076GAT(2340) ; 6076GAT(2340)*
g4700 not 6073GAT(2341) ; 6073GAT(2341)*
g4701 not 6070GAT(2342) ; 6070GAT(2342)*
g4702 not 6068GAT(2343) ; 6068GAT(2343)*
g4703 not 6069GAT(2345) ; 6069GAT(2345)*
g4704 not 6064GAT(2346) ; 6064GAT(2346)*
g4705 not 6061GAT(2344) ; 6061GAT(2344)*
g4706 not 588GAT(272) ; 588GAT(272)*
g4707 not 6101GAT(2348) ; 6101GAT(2348)*
g4708 not 6102GAT(2349) ; 6102GAT(2349)*
g4709 not 6097GAT(2350) ; 6097GAT(2350)*
g4710 not 6094GAT(2351) ; 6094GAT(2351)*
g4711 not 6091GAT(2352) ; 6091GAT(2352)*
g4712 not 6089GAT(2353) ; 6089GAT(2353)*
g4713 not 6090GAT(2354) ; 6090GAT(2354)*
g4714 not 6085GAT(2355) ; 6085GAT(2355)*
g4715 not 6118GAT(2357) ; 6118GAT(2357)*
g4716 not 6119GAT(2358) ; 6119GAT(2358)*
g4717 not 6114GAT(2359) ; 6114GAT(2359)*
g4718 not 6111GAT(2360) ; 6111GAT(2360)*
g4719 not 6108GAT(2362) ; 6108GAT(2362)*
g4720 not 6106GAT(2361) ; 6106GAT(2361)*
g4721 not 6107GAT(2363) ; 6107GAT(2363)*
g4722 not 6128GAT(2365) ; 6128GAT(2365)*
g4723 not 6129GAT(2366) ; 6129GAT(2366)*
g4724 not 6124GAT(2367) ; 6124GAT(2367)*
g4725 not 6133GAT(2370) ; 6133GAT(2370)*
g4726 not 6134GAT(2371) ; 6134GAT(2371)*
g4727 not 6141GAT(2373) ; 6141GAT(2373)*
g4728 not 6138GAT(2372) ; 6138GAT(2372)*
g4729 not 6135GAT(2369) ; 6135GAT(2369)*
g4730 not 6147GAT(2374) ; 6147GAT(2374)*
g4731 not 6145GAT(2375) ; 6145GAT(2375)*
g4732 not 6146GAT(2376) ; 6146GAT(2376)*
g4733 not 6151GAT(2377) ; 6151GAT(2377)*
g4734 not 6130GAT(2364) ; 6130GAT(2364)*
g4735 not 6157GAT(2379) ; 6157GAT(2379)*
g4736 not 6155GAT(2380) ; 6155GAT(2380)*
g4737 not 6156GAT(2381) ; 6156GAT(2381)*
g4738 not 6161GAT(2382) ; 6161GAT(2382)*
g4739 not 6120GAT(2356) ; 6120GAT(2356)*
g4740 not 6167GAT(2384) ; 6167GAT(2384)*
g4741 not 6165GAT(2385) ; 6165GAT(2385)*
g4742 not 6166GAT(2386) ; 6166GAT(2386)*
g4743 not 6171GAT(2387) ; 6171GAT(2387)*
g4744 not 6103GAT(2347) ; 6103GAT(2347)*
g4745 not 6177GAT(2389) ; 6177GAT(2389)*
g4746 not 6175GAT(2390) ; 6175GAT(2390)*
g4747 not 6176GAT(2391) ; 6176GAT(2391)*
g4748 not 6181GAT(2392) ; 6181GAT(2392)*
g4749 not 6082GAT(2337) ; 6082GAT(2337)*
g4750 not 6187GAT(2394) ; 6187GAT(2394)*
g4751 not 6185GAT(2395) ; 6185GAT(2395)*
g4752 not 6186GAT(2396) ; 6186GAT(2396)*
g4753 not 6191GAT(2397) ; 6191GAT(2397)*
g4754 not 6058GAT(2325) ; 6058GAT(2325)*
g4755 not 6197GAT(2399) ; 6197GAT(2399)*
g4756 not 6195GAT(2400) ; 6195GAT(2400)*
g4757 not 6196GAT(2401) ; 6196GAT(2401)*
g4758 not 6201GAT(2402) ; 6201GAT(2402)*
g4759 not 6032GAT(2312) ; 6032GAT(2312)*
g4760 not 6207GAT(2404) ; 6207GAT(2404)*
g4761 not 6205GAT(2405) ; 6205GAT(2405)*
g4762 not 6206GAT(2406) ; 6206GAT(2406)*
g4763 not 6211GAT(2407) ; 6211GAT(2407)*
g4764 not 6002GAT(2297) ; 6002GAT(2297)*
g4765 not 6217GAT(2409) ; 6217GAT(2409)*
g4766 not 6215GAT(2410) ; 6215GAT(2410)*
g4767 not 6216GAT(2411) ; 6216GAT(2411)*
g4768 not 6221GAT(2412) ; 6221GAT(2412)*
g4769 not 5968GAT(2277) ; 5968GAT(2277)*
g4770 not 6227GAT(2414) ; 6227GAT(2414)*
g4771 not 6225GAT(2415) ; 6225GAT(2415)*
g4772 not 6226GAT(2416) ; 6226GAT(2416)*
g4773 not 6231GAT(2417) ; 6231GAT(2417)*
g4774 not 5925GAT(2258) ; 5925GAT(2258)*
g4775 not 6237GAT(2419) ; 6237GAT(2419)*
g4776 not 6235GAT(2420) ; 6235GAT(2420)*
g4777 not 6236GAT(2421) ; 6236GAT(2421)*
g4778 not 6241GAT(2422) ; 6241GAT(2422)*
g4779 not 5879GAT(2238) ; 5879GAT(2238)*
g4780 not 6247GAT(2424) ; 6247GAT(2424)*
g4781 not 6245GAT(2425) ; 6245GAT(2425)*
g4782 not 6246GAT(2426) ; 6246GAT(2426)*
g4783 not 6251GAT(2427) ; 6251GAT(2427)*
g4784 not 5831GAT(2215) ; 5831GAT(2215)*
g4785 not 6257GAT(2429) ; 6257GAT(2429)*
g4786 not 6255GAT(2430) ; 6255GAT(2430)*
g4787 not 6256GAT(2431) ; 6256GAT(2431)*
g4788 not 6261GAT(2432) ; 6261GAT(2432)*
g4789 not 5782GAT(2192) ; 5782GAT(2192)*
g4790 not 6267GAT(2434) ; 6267GAT(2434)*
g4791 not 6265GAT(2435) ; 6265GAT(2435)*
g4792 not 6266GAT(2436) ; 6266GAT(2436)*
g4793 not 6271GAT(2437) ; 6271GAT(2437)*
g4794 not 5727GAT(2167) ; 5727GAT(2167)*
g4795 not 6277GAT(2439) ; 6277GAT(2439)*
g4796 not 6275GAT(2440) ; 6275GAT(2440)*
g4797 not 6276GAT(2441) ; 6276GAT(2441)*
g4798 not 6281GAT(2442) ; 6281GAT(2442)*
g4799 not 6285GAT(2445) ; 6285GAT(2445)*
g4800 not 6286GAT(2446) ; 6286GAT(2446)*
