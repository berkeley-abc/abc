name C2670.iscas
i 1(0)
i 2(1)
i 3(2)
i 4(3)
i 5(4)
i 6(5)
i 7(6)
i 8(7)
i 11(8)
i 14(9)
i 15(10)
i 16(11)
i 19(12)
i 20(13)
i 21(14)
i 22(15)
i 23(16)
i 24(17)
i 25(18)
i 26(19)
i 27(20)
i 28(21)
i 29(22)
i 32(23)
i 33(24)
i 34(25)
i 35(26)
i 36(27)
i 37(28)
i 40(29)
i 43(30)
i 44(31)
i 47(32)
i 48(33)
i 49(34)
i 50(35)
i 51(36)
i 52(37)
i 53(38)
i 54(39)
i 55(40)
i 56(41)
i 57(42)
i 60(43)
i 61(44)
i 62(45)
i 63(46)
i 64(47)
i 65(48)
i 66(49)
i 67(50)
i 68(51)
i 69(52)
i 72(53)
i 73(54)
i 74(55)
i 75(56)
i 76(57)
i 77(58)
i 78(59)
i 79(60)
i 80(61)
i 81(62)
i 82(63)
i 85(64)
i 86(65)
i 87(66)
i 88(67)
i 89(68)
i 90(69)
i 91(70)
i 92(71)
i 93(72)
i 94(73)
i 95(74)
i 96(75)
i 99(76)
i 100(77)
i 101(78)
i 102(79)
i 103(80)
i 104(81)
i 105(82)
i 106(83)
i 107(84)
i 108(85)
i 111(86)
i 112(87)
i 113(88)
i 114(89)
i 115(90)
i 116(91)
i 117(92)
i 118(93)
i 119(94)
i 120(95)
i 123(96)
i 124(97)
i 125(98)
i 126(99)
i 127(100)
i 128(101)
i 129(102)
i 130(103)
i 131(104)
i 132(105)
i 135(106)
i 136(107)
i 137(108)
i 138(109)
i 139(110)
i 140(111)
i 141(112)
i 142(113)
i IN-169(114)
i IN-174(115)
i IN-177(116)
i IN-178(117)
i IN-179(118)
i IN-180(119)
i IN-181(120)
i IN-182(121)
i IN-183(122)
i IN-184(123)
i IN-185(124)
i IN-186(125)
i IN-189(126)
i IN-190(127)
i IN-191(128)
i IN-192(129)
i IN-193(130)
i IN-194(131)
i IN-195(132)
i IN-196(133)
i IN-197(134)
i IN-198(135)
i IN-199(136)
i IN-200(137)
i IN-201(138)
i IN-202(139)
i IN-203(140)
i IN-204(141)
i IN-205(142)
i IN-206(143)
i IN-207(144)
i IN-208(145)
i IN-209(146)
i IN-210(147)
i IN-211(148)
i IN-212(149)
i IN-213(150)
i IN-214(151)
i IN-215(152)
i IN-239(153)
i IN-240(154)
i IN-241(155)
i IN-242(156)
i IN-243(157)
i IN-244(158)
i IN-245(159)
i IN-246(160)
i IN-247(161)
i IN-248(162)
i IN-249(163)
i IN-250(164)
i IN-251(165)
i IN-252(166)
i IN-253(167)
i IN-254(168)
i IN-255(169)
i IN-256(170)
i IN-257(171)
i IN-262(172)
i IN-263(173)
i IN-264(174)
i IN-265(175)
i IN-266(176)
i IN-267(177)
i IN-268(178)
i IN-269(179)
i IN-270(180)
i IN-271(181)
i IN-272(182)
i IN-273(183)
i IN-274(184)
i IN-275(185)
i IN-276(186)
i IN-277(187)
i IN-278(188)
i IN-279(189)
i 452(190)
i 483(191)
i 543(192)
i 559(193)
i 567(194)
i 651(195)
i 661(196)
i 860(197)
i 868(198)
i 1083(199)
i 1341(200)
i 1348(201)
i 1384(202)
i 1956(203)
i 1961(204)
i 1966(205)
i 1971(206)
i 1976(207)
i 1981(208)
i 1986(209)
i 1991(210)
i 1996(211)
i 2066(212)
i 2067(213)
i 2072(214)
i 2078(215)
i 2084(216)
i 2090(217)
i 2096(218)
i 2100(219)
i 2104(220)
i 2105(221)
i 2106(222)
i 2427(223)
i 2430(224)
i 2435(225)
i 2438(226)
i 2443(227)
i 2446(228)
i 2451(229)
i 2454(230)
i 2474(231)
i 2678(232)

o 169(114)
o 174(115)
o 177(116)
o 178(117)
o 179(118)
o 180(119)
o 181(120)
o 182(121)
o 183(122)
o 184(123)
o 185(124)
o 186(125)
o 189(126)
o 190(127)
o 191(128)
o 192(129)
o 193(130)
o 194(131)
o 195(132)
o 196(133)
o 197(134)
o 198(135)
o 199(136)
o 200(137)
o 201(138)
o 202(139)
o 203(140)
o 204(141)
o 205(142)
o 206(143)
o 207(144)
o 208(145)
o 209(146)
o 210(147)
o 211(148)
o 212(149)
o 213(150)
o 214(151)
o 215(152)
o 239(153)
o 240(154)
o 241(155)
o 242(156)
o 243(157)
o 244(158)
o 245(159)
o 246(160)
o 247(161)
o 248(162)
o 249(163)
o 250(164)
o 251(165)
o 252(166)
o 253(167)
o 254(168)
o 255(169)
o 256(170)
o 257(171)
o 262(172)
o 263(173)
o 264(174)
o 265(175)
o 266(176)
o 267(177)
o 268(178)
o 269(179)
o 270(180)
o 271(181)
o 272(182)
o 273(183)
o 274(184)
o 275(185)
o 276(186)
o 277(187)
o 278(188)
o 279(189)
o 350(301)
o 335(299)
o 409(298)
o 369(289)
o 367(288)
o 411(264)
o 337(263)
o 384(262)
o 218(311)
o 219(302)
o 220(306)
o 221(305)
o 235(307)
o 236(303)
o 237(309)
o 238(304)
o 158(349)
o 259(414)
o 391(379)
o 173(389)
o 223(413)
o 234(376)
o 217(423)
o 325(507)
o 261(506)
o 319(656)
o 160(609)
o 162(612)
o 164(607)
o 166(625)
o 168(623)
o 171(621)
o 153(671)
o 176(803)
o 188(761)
o 299(692)
o 301(694)
o 286(696)
o 303(698)
o 288(700)
o 305(702)
o 290(704)
o 284(847)
o 321(848)
o 297(849)
o 280(850)
o 148(851)
o 282(922)
o 323(923)
o 156(1046)
o 401(1276)
o 227(1179)
o 229(1180)
o 311(1278)
o 150(1277)
o 145(1358)
o 395(1392)
o 295(1400)
o 331(1401)
o 397(1406)
o 329(1414)
o 231(1422)
o 308(1425)
o 225(1424)

g1 not 44(31) ; 218(311)
g2 not 132(105) ; 219(302)
g3 not 82(63) ; 220(306)
g4 not 96(75) ; 221(305)
g5 not 69(52) ; 235(307)
g6 not 120(95) ; 236(303)
g7 not 57(42) ; 237(309)
g8 not 108(85) ; 238(304)
g9 not 157(259) ; 158(349)
g10 not 258(321) ; 259(414)
g11 and 391(379) 94(73) ; 173(389)
g12 not 1955(320) ; 223(413)
g13 or 1955(320)* 567(194)* ; 234(376)
g14 not 216(333) ; 217(423)
g15 not 325(507) ; 261(506)
g16 not 1464(560) ; 160(609)
g17 not 1467(561) ; 162(612)
g18 not 1461(559) ; 164(607)
g19 not 1329(569) ; 166(625)
g20 not 1327(568) ; 168(623)
g21 not 857(567) ; 171(621)
g22 or 152(599) 865(291) ; 153(671)
g23 not 175(710) ; 176(803)
g24 not 187(673) ; 188(761)
g25 or 147(600) 146(758) ; 148(851)
g26 or 155(967)* 154(964)* ; 156(1046)
g27 not 1830(1108) ; 227(1179)
g28 not 1553(1110) ; 229(1180)
g29 not 311(1278) ; 150(1277)
g30 or 144(601) 143(1330) ; 145(1358)
g31 not 473(1420) ; 231(1422)
g32 not 308(1425) ; 225(1424)
g33 not 2678(232) ; 2682(233)
g34 not 2474(231) ; 2478(234)
g35 not 2454(230) ; 2458(235)
g36 not 2451(229) ; 2457(236)
g37 not 2446(228) ; 2450(237)
g38 not 2443(227) ; 2449(238)
g39 not 2438(226) ; 2442(239)
g40 not 2435(225) ; 2441(240)
g41 not 2430(224) ; 2434(241)
g42 not 2427(223) ; 2433(242)
g43 and 2105(221) ; 1655(243)
g44 and 2105(221) ; 1418(244)
g45 and 2104(220) ; 1631(245)
g46 and 2104(220) ; 1394(246)
g47 not 2100(219) ; 2103(247)
g48 and 2100(219) ; 2699(248)
g49 not 2096(218) ; 2099(249)
g50 and 2096(218) ; 2702(250)
g51 not 2090(217) ; 2094(251)
g52 and 2090(217) ; 2691(252)
g53 not 2084(216) ; 2088(253)
g54 and 2084(216) ; 2694(254)
g55 not 2078(215) ; 2082(255)
g56 and 2078(215) ; 2683(256)
g57 not 2072(214) ; 2076(257)
g58 and 2072(214) ; 2686(258)
g59 and 2072(214) 2078(215) 2084(216) 2090(217) ; 157(259)
g60 not 2067(213) ; 2070(260)
g61 and 2067(213) ; 2675(261)
g62 not 1996(211) ; 1999(265)
g63 and 1996(211) ; 2505(266)
g64 not 1991(210) ; 1994(267)
g65 and 1991(210) ; 2508(268)
g66 not 1986(209) ; 1989(269)
g67 and 1986(209) ; 2495(270)
g68 not 1981(208) ; 1984(271)
g69 and 1981(208) ; 2498(272)
g70 not 1976(207) ; 1979(273)
g71 and 1976(207) ; 2487(274)
g72 not 1971(206) ; 1974(275)
g73 and 1971(206) ; 2490(276)
g74 not 1966(205) ; 1969(277)
g75 and 1966(205) ; 2479(278)
g76 not 1961(204) ; 1964(279)
g77 and 1961(204) ; 2482(280)
g78 not 1956(203) ; 1959(281)
g79 and 1956(203) ; 2471(282)
g80 not 1384(202) ; 1385(283)
g81 not 1348(201) ; 1351(284)
g82 and 1348(201) ; 2461(285)
g83 not 1341(200) ; 1344(286)
g84 and 1341(200) ; 2464(287)
g85 not 868(198) ; 875(290)
g86 not 860(197) ; 865(291)
g87 and 661(196) ; 480(292)
g88 and 651(195) ; 1284(293)
g89 and 651(195) ; 795(294)
g90 not 559(193) ; 560(295)
g91 and 543(192) ; 1261(296)
g92 and 543(192) ; 772(297)
g93 and 452(190) ; 391(379)
g94 and 69(52) 108(85) 57(42) 120(95) ; 1254(308)
g95 and 44(31) 96(75) 82(63) 132(105) ; 1251(310)
g96 and 37(28) ; 486(312)
g97 and 29(22) ; 2012(313)
g98 and 29(22) ; 2001(314)
g99 and 16(11) ; 1721(315)
g100 and 16(11) ; 1710(316)
g101 and 868(198) 11(8) ; 882(317)
g102 and 8(7) ; 658(318)
g103 and 8(7) ; 655(319)
g104 and 661(196) 7(6) ; 1955(320)
g105 and 661(196) 15(10) 2(1) ; 258(321)
g106 and 3(2) 1(0) ; 546(322)
g107 or 2682(233)* 2675(261)* ; 1776(323)
g108 or 2478(234)* 2471(282)* ; 1499(324)
g109 or 2457(236)* 2454(230)* ; 2459(325)
g110 or 2458(235)* 2451(229)* ; 2460(326)
g111 or 2449(238)* 2446(228)* ; 1493(327)
g112 or 2450(237)* 2443(227)* ; 1494(328)
g113 or 2441(240)* 2438(226)* ; 1484(329)
g114 or 2442(239)* 2435(225)* ; 1485(330)
g115 or 2433(242)* 2430(224)* ; 1475(331)
g116 or 2434(241)* 2427(223)* ; 1476(332)
g117 and 1955(320) 2106(222) ; 216(333)
g118 not 1655(243) ; 1667(334)
g119 and 1418(244) 1394(246) ; 1460(335)
g120 not 1418(244) ; 1430(336)
g121 not 1631(245) ; 1643(337)
g122 not 1394(246) ; 1406(338)
g123 not 2699(248) ; 2705(339)
g124 not 2702(250) ; 2706(340)
g125 and 2094(251) ; 2775(341)
g126 not 2691(252) ; 2697(342)
g127 and 2088(253) ; 2767(343)
g128 not 2694(254) ; 2698(344)
g129 and 2082(255) ; 2759(345)
g130 not 2683(256) ; 2689(346)
g131 and 2076(257) ; 2751(347)
g132 not 2686(258) ; 2690(348)
g133 and 2070(260) ; 2743(350)
g134 not 2675(261) ; 2681(351)
g135 and 1999(265) ; 2735(352)
g136 not 2505(266) ; 2511(353)
g137 and 1994(267) ; 2623(354)
g138 not 2508(268) ; 2512(355)
g139 and 1989(269) ; 2615(356)
g140 not 2495(270) ; 2501(357)
g141 and 1984(271) ; 2607(358)
g142 not 2498(272) ; 2502(359)
g143 and 1979(273) ; 2599(360)
g144 not 2487(274) ; 2493(361)
g145 and 1974(275) ; 2591(362)
g146 not 2490(276) ; 2494(363)
g147 and 1969(277) ; 2583(364)
g148 not 2479(278) ; 2485(365)
g149 and 1964(279) ; 2575(366)
g150 not 2482(280) ; 2486(367)
g151 and 1959(281) ; 2567(368)
g152 not 2471(282) ; 2477(369)
g153 and 1351(284) ; 2559(370)
g154 not 2461(285) ; 2467(371)
g155 and 1344(286) ; 2551(372)
g156 not 2464(287) ; 2468(373)
g157 not 1284(293) ; 1296(374)
g158 not 795(294) ; 807(375)
g159 not 1261(296) ; 1273(377)
g160 not 772(297) ; 784(378)
g161 and 1655(243) 1631(245) 118(93) ; 1681(380)
g162 and 1655(243) 1631(245) 117(92) ; 1689(381)
g163 and 1655(243) 1631(245) 116(91) ; 1693(382)
g164 and 1655(243) 1631(245) 115(90) ; 1697(383)
g165 and 1418(244) 1394(246) 114(89) ; 1444(384)
g166 and 1418(244) 1394(246) 113(88) ; 1448(385)
g167 and 1418(244) 1394(246) 112(87) ; 1452(386)
g168 and 1418(244) 1394(246) 111(86) ; 1456(387)
g169 and 1655(243) 1631(245) 107(84) ; 1685(388)
g170 and 795(294) 772(297) 80(61) ; 821(390)
g171 and 795(294) 772(297) 79(60) ; 829(391)
g172 and 795(294) 772(297) 78(59) ; 833(392)
g173 and 795(294) 772(297) 77(58) ; 837(393)
g174 and 1284(293) 1261(296) 76(57) ; 1310(394)
g175 and 1284(293) 1261(296) 75(56) ; 1314(395)
g176 and 1284(293) 1261(296) 74(55) ; 1318(396)
g177 and 1284(293) 1261(296) 73(54) ; 1322(397)
g178 and 1284(293) 1261(296) 72(53) ; 1326(398)
g179 and 795(294) 772(297) 68(51) ; 825(399)
g180 and 1251(310) 1254(308) ; 325(507)
g181 not 1254(308) ; 1256(401)
g182 not 1251(310) ; 1253(402)
g183 not 486(312) ; 487(403)
g184 not 2012(313) ; 2018(404)
g185 not 2001(314) ; 2007(405)
g186 not 1721(315) ; 1728(406)
g187 not 1710(316) ; 1716(407)
g188 and 875(290) 11(8) ; 881(408)
g189 and 658(318) ; 1831(409)
g190 and 658(318) ; 1893(410)
g191 and 655(319) ; 748(411)
g192 and 655(319) ; 994(412)
g193 not 546(322) ; 547(415)
g194 or 2681(351)* 2678(232)* ; 1775(416)
g195 or 2477(369)* 2474(231)* ; 1498(417)
g196 or 2460(326)* 2459(325)* ; 2518(418)
g197 or 1494(328)* 1493(327)* ; 1495(419)
g198 or 1485(330)* 1484(329)* ; 1486(420)
g199 or 1476(332)* 1475(331)* ; 1477(421)
g200 and 1253(402) 2106(222) ; 550(422)
g201 and 1418(244) 1406(338) ; 1459(424)
g202 and 1430(336) 1406(338) ; 1457(425)
g203 and 1430(336) 1394(246) ; 1458(426)
g204 or 2706(340)* 2699(248)* ; 2708(427)
g205 or 2705(339)* 2702(250)* ; 2707(428)
g206 not 2775(341) ; 2781(429)
g207 or 2698(344)* 2691(252)* ; 1794(430)
g208 not 2767(343) ; 2773(431)
g209 or 2697(342)* 2694(254)* ; 1793(432)
g210 not 2759(345) ; 2765(433)
g211 or 2690(348)* 2683(256)* ; 1785(434)
g212 not 2751(347) ; 2757(435)
g213 or 2689(346)* 2686(258)* ; 1784(436)
g214 not 2743(350) ; 2749(437)
g215 not 2735(352) ; 2741(438)
g216 or 2512(355)* 2505(266)* ; 2514(439)
g217 not 2623(354) ; 2629(440)
g218 or 2511(353)* 2508(268)* ; 2513(441)
g219 not 2615(356) ; 2621(442)
g220 or 2502(359)* 2495(270)* ; 2504(443)
g221 not 2607(358) ; 2613(444)
g222 or 2501(357)* 2498(272)* ; 2503(445)
g223 not 2599(360) ; 2605(446)
g224 or 2494(363)* 2487(274)* ; 1517(447)
g225 not 2591(362) ; 2597(448)
g226 or 2493(361)* 2490(276)* ; 1516(449)
g227 not 2583(364) ; 2589(450)
g228 or 2486(367)* 2479(278)* ; 1508(451)
g229 not 2575(366) ; 2581(452)
g230 or 2485(365)* 2482(280)* ; 1507(453)
g231 not 2567(368) ; 2573(454)
g232 not 2559(370) ; 2565(455)
g233 or 2468(373)* 2461(285)* ; 2470(456)
g234 not 2551(372) ; 2557(457)
g235 or 2467(371)* 2464(287)* ; 2469(458)
g236 and 1284(293) 1273(377) ; 1317(459)
g237 and 1256(401) 567(194) ; 552(460)
g238 and 1667(334) 1643(337) 142(113) ; 1678(461)
g239 and 1667(334) 1643(337) 141(112) ; 1686(462)
g240 and 1667(334) 1643(337) 140(111) ; 1690(463)
g241 and 1667(334) 1643(337) 139(110) ; 1694(464)
g242 and 1430(336) 1406(338) 138(109) ; 1441(465)
g243 and 1430(336) 1406(338) 137(108) ; 1445(466)
g244 and 1430(336) 1406(338) 136(107) ; 1449(467)
g245 and 1430(336) 1406(338) 135(106) ; 1453(468)
g246 and 1667(334) 1643(337) 131(104) ; 1682(469)
g247 and 1655(243) 1643(337) 130(103) ; 1680(470)
g248 and 1655(243) 1643(337) 129(102) ; 1688(471)
g249 and 1655(243) 1643(337) 128(101) ; 1692(472)
g250 and 1655(243) 1643(337) 127(100) ; 1696(473)
g251 and 1418(244) 1406(338) 126(99) ; 1443(474)
g252 and 1418(244) 1406(338) 125(98) ; 1447(475)
g253 and 1418(244) 1406(338) 124(97) ; 1451(476)
g254 and 1418(244) 1406(338) 123(96) ; 1455(477)
g255 and 1655(243) 1643(337) 119(94) ; 1684(478)
g256 and 1667(334) 1631(245) 106(83) ; 1679(479)
g257 and 1667(334) 1631(245) 105(82) ; 1687(480)
g258 and 1667(334) 1631(245) 104(81) ; 1691(481)
g259 and 1667(334) 1631(245) 103(80) ; 1695(482)
g260 and 1430(336) 1394(246) 102(79) ; 1442(483)
g261 and 1430(336) 1394(246) 101(78) ; 1446(484)
g262 and 1430(336) 1394(246) 100(77) ; 1450(485)
g263 and 1430(336) 1394(246) 99(76) ; 1454(486)
g264 and 1667(334) 1631(245) 95(74) ; 1683(487)
g265 and 807(375) 784(378) 93(72) ; 818(488)
g266 and 807(375) 784(378) 92(71) ; 826(489)
g267 and 807(375) 784(378) 91(70) ; 830(490)
g268 and 807(375) 784(378) 90(69) ; 834(491)
g269 and 1296(374) 1273(377) 89(68) ; 1307(492)
g270 and 1296(374) 1273(377) 88(67) ; 1311(493)
g271 and 1296(374) 1273(377) 87(66) ; 1315(494)
g272 and 1296(374) 1273(377) 86(65) ; 1319(495)
g273 and 1296(374) 1273(377) 85(64) ; 1323(496)
g274 and 807(375) 784(378) 81(62) ; 822(497)
g275 and 795(294) 784(378) 67(50) ; 820(498)
g276 and 795(294) 784(378) 66(49) ; 828(499)
g277 and 795(294) 784(378) 65(48) ; 832(500)
g278 and 795(294) 784(378) 64(47) ; 836(501)
g279 and 1284(293) 1273(377) 63(46) ; 1309(502)
g280 and 1284(293) 1273(377) 62(45) ; 1313(503)
g281 and 1284(293) 1273(377) 61(44) ; 1321(504)
g282 and 1284(293) 1273(377) 60(43) ; 1325(505)
g283 and 795(294) 784(378) 56(41) ; 824(508)
g284 and 807(375) 772(297) 55(40) ; 819(509)
g285 and 807(375) 772(297) 54(39) ; 827(510)
g286 and 807(375) 772(297) 53(38) ; 831(511)
g287 and 807(375) 772(297) 52(37) ; 835(512)
g288 and 1296(374) 1261(296) 51(36) ; 1308(513)
g289 and 1296(374) 1261(296) 50(35) ; 1312(514)
g290 and 1296(374) 1261(296) 49(34) ; 1316(515)
g291 and 1296(374) 1261(296) 48(33) ; 1320(516)
g292 and 1296(374) 1261(296) 47(32) ; 1324(517)
g293 and 807(375) 772(297) 43(30) ; 823(518)
g294 and 2018(404) 35(26) ; 2035(519)
g295 and 2018(404) 34(25) ; 2033(520)
g296 and 2007(405) 33(24) ; 2029(521)
g297 and 2007(405) 32(23) ; 2025(522)
g298 and 2018(404) 28(21) ; 2037(523)
g299 and 2018(404) 27(20) ; 2031(524)
g300 and 2007(405) 26(19) ; 2027(525)
g301 and 2007(405) 25(18) ; 2023(526)
g302 and 1728(406) 24(17) ; 1750(527)
g303 and 1728(406) 23(16) ; 1746(528)
g304 and 1728(406) 22(15) ; 1744(529)
g305 and 1728(406) 21(14) ; 1742(530)
g306 and 1716(407) 20(13) ; 1738(531)
g307 and 1716(407) 19(12) ; 1734(532)
g308 or 882(317) 881(408) ; 894(533)
g309 and 1728(406) 6(5) ; 1748(534)
g310 and 1716(407) 5(4) ; 1740(535)
g311 and 1716(407) 4(3) ; 1736(536)
g312 or 1776(323)* 1775(416)* ; 1777(537)
g313 or 1499(324)* 1498(417)* ; 1500(538)
g314 not 2518(418) ; 2522(539)
g315 and 1495(419) ; 1525(540)
g316 and 1495(419) ; 1521(541)
g317 not 1486(420) ; 1490(542)
g318 not 1477(421) ; 1481(543)
g319 not 550(422) ; 551(544)
g320 or 1460(335) 1459(424) 1458(426) 1457(425) ; 1473(545)
g321 or 2708(427)* 2707(428)* ; 2730(546)
g322 or 1794(430)* 1793(432)* ; 1795(547)
g323 or 1785(434)* 1784(436)* ; 1786(548)
g324 or 2514(439)* 2513(441)* ; 2525(549)
g325 or 2504(443)* 2503(445)* ; 2528(550)
g326 or 1517(447)* 1516(449)* ; 1518(551)
g327 or 1508(451)* 1507(453)* ; 1509(552)
g328 or 2470(456)* 2469(458)* ; 2515(553)
g329 not 552(460) ; 553(554)
g330 or 1681(380) 1680(470) 1679(479) 1678(461) ; 2634(555)
g331 or 1689(381) 1688(471) 1687(480) 1686(462) ; 1701(556)
g332 or 1693(382) 1692(472) 1691(481) 1690(463) ; 1704(557)
g333 or 1697(383) 1696(473) 1695(482) 1694(464) ; 1707(558)
g334 or 1444(384) 1443(474) 1442(483) 1441(465) ; 1461(559)
g335 or 1448(385) 1447(475) 1446(484) 1445(466) ; 1464(560)
g336 or 1452(386) 1451(476) 1450(485) 1449(467) ; 1467(561)
g337 or 1456(387) 1455(477) 1454(486) 1453(468) ; 1470(562)
g338 or 1685(388) 1684(478) 1683(487) 1682(469) ; 1698(563)
g339 or 821(390) 820(498) 819(509) 818(488) ; 838(564)
g340 or 829(391) 828(499) 827(510) 826(489) ; 846(565)
g341 or 833(392) 832(500) 831(511) 830(490) ; 854(566)
g342 or 837(393) 836(501) 835(512) 834(491) ; 857(567)
g343 or 1310(394) 1309(502) 1308(513) 1307(492) ; 1327(568)
g344 or 1314(395) 1313(503) 1312(514) 1311(493) ; 1329(569)
g345 or 1318(396) 1317(459) 1316(515) 1315(494) ; 1331(570)
g346 or 1322(397) 1321(504) 1320(516) 1319(495) ; 1333(571)
g347 or 1326(398) 1325(505) 1324(517) 1323(496) ; 1335(572)
g348 or 825(399) 824(508) 823(518) 822(497) ; 841(573)
g349 not 1777(537) ; 1781(574)
g350 not 1500(538) ; 1504(575)
g351 or 2522(539)* 2515(553)* ; 2524(576)
g352 and 1525(540) 1481(543) 1490(542) ; 1541(577)
g353 not 1525(540) ; 1528(578)
g354 not 1521(541) ; 1524(579)
g355 and 1521(541) 1477(421) 1486(420) ; 1538(580)
g356 and 553(554) 551(544) ; 319(656)
g357 and 1473(545) ; 2665(582)
g358 or 1473(545)* 2103(247)* ; 1218(583)
g359 not 2730(546) ; 2734(584)
g360 or 1470(562)* 2099(249)* ; 1213(585)
g361 and 1795(547) ; 1810(586)
g362 and 1795(547) ; 1806(587)
g363 not 1786(548) ; 1790(588)
g364 not 2525(549) ; 2531(589)
g365 not 2528(550) ; 2532(590)
g366 and 1518(551) ; 1533(591)
g367 and 1518(551) ; 1529(592)
g368 not 1509(552) ; 1513(593)
g369 and 1385(283) 1461(559) ; 1387(594)
g370 not 2515(553) ; 2521(595)
g371 and 875(290) 841(573) ; 885(596)
g372 and 875(290) 846(565) ; 887(597)
g373 and 868(198) 1327(568) ; 893(598)
g374 and 860(197) 841(573) ; 152(599)
g375 and 860(197) 846(565) ; 147(600)
g376 and 860(197) 838(564) ; 144(601)
g377 not 2634(555) ; 2638(602)
g378 and 1701(556) ; 2642(603)
g379 and 1704(557) ; 1250(604)
g380 and 1704(557) ; 2639(605)
g381 and 1707(558) ; 2650(606)
g382 and 1461(559) ; 2647(608)
g383 not 1464(560) ; 1389(610)
g384 and 1464(560) ; 2658(611)
g385 and 1467(561) ; 2655(613)
g386 and 1470(562) ; 2668(614)
g387 and 1698(563) ; 2631(615)
g388 and 838(564) ; 516(616)
g389 not 838(564) ; 1028(617)
g390 not 846(565) ; 1035(618)
g391 not 846(565) ; 852(619)
g392 and 854(566) ; 299(692)
g393 and 857(567) ; 301(694)
g394 and 1327(568) ; 286(696)
g395 and 1329(569) ; 303(698)
g396 and 1331(570) ; 288(700)
g397 and 1333(571) ; 305(702)
g398 and 1335(572) ; 290(704)
g399 not 841(573) ; 1031(630)
g400 and 841(573) ; 2154(631)
g401 and 2012(313) 1467(561) ; 2036(632)
g402 and 2012(313) 1464(560) ; 2034(633)
g403 and 2012(313) 1461(559) ; 2032(634)
g404 and 2012(313) 1470(562) ; 2038(635)
g405 and 2001(314) 1698(563) ; 2024(636)
g406 and 2001(314) 1707(558) ; 2030(637)
g407 and 2001(314) 1704(557) ; 2028(638)
g408 and 2001(314) 1701(556) ; 2026(639)
g409 and 1721(315) 1331(570) ; 1747(640)
g410 and 1721(315) 1329(569) ; 1745(641)
g411 and 1721(315) 1327(568) ; 1743(642)
g412 and 1721(315) 1335(572) ; 1751(643)
g413 and 1721(315) 1333(571) ; 1749(644)
g414 and 1710(316) 841(573) ; 1735(645)
g415 and 1710(316) 857(567) ; 1741(646)
g416 and 1710(316) 854(566) ; 1739(647)
g417 and 1710(316) 846(565) ; 1737(648)
g418 and 1806(587) 1777(537) 1786(548) ; 1821(649)
g419 and 1810(586) 1781(574) 1790(588) ; 1824(650)
g420 and 1529(592) 1500(538) 1509(552) ; 1544(651)
g421 and 1533(591) 1504(575) 1513(593) ; 1547(652)
g422 or 2521(595)* 2518(418)* ; 2523(653)
g423 and 1524(579) 1486(420) 1481(543) ; 1537(654)
g424 and 1528(578) 1490(542) 1477(421) ; 1540(655)
g425 and 1473(545) 1218(583) ; 1234(657)
g426 not 2665(582) ; 2671(658)
g427 and 1218(583) 2103(247) ; 1232(659)
g428 and 1213(585) 2099(249) ; 1225(660)
g429 not 1810(586) ; 1813(661)
g430 not 1806(587) ; 1809(662)
g431 or 2532(590)* 2525(549)* ; 2534(663)
g432 or 2531(589)* 2528(550)* ; 2533(664)
g433 not 1533(591) ; 1536(665)
g434 not 1529(592) ; 1532(666)
g435 not 1387(594) ; 466(667)
g436 and 875(290) 516(616) ; 883(668)
g437 and 875(290) 299(692) ; 891(669)
g438 and 868(198) 301(694) ; 889(670)
g439 or 852(619)* 560(295)* ; 562(672)
g440 and 547(415) 319(656) 483(191) 480(292) ; 187(673)
g441 or 2638(602)* 2631(615)* ; 1753(674)
g442 not 2642(603) ; 2646(675)
g443 not 2639(605) ; 2645(676)
g444 not 2650(606) ; 2654(677)
g445 not 2647(608) ; 2653(678)
g446 not 2658(611) ; 2662(679)
g447 not 2655(613) ; 2661(680)
g448 and 1470(562) 1213(585) ; 1227(681)
g449 not 2668(614) ; 2672(682)
g450 not 2631(615) ; 2637(683)
g451 and 516(616) ; 2235(684)
g452 and 1028(617) ; 2110(685)
g453 and 1028(617) ; 2164(686)
g454 and 1035(618) ; 2350(687)
g455 and 1035(618) ; 2118(688)
g456 and 1035(618) ; 2262(689)
g457 and 1035(618) ; 2172(690)
g458 not 852(619) ; 2151(691)
g459 not 299(692) ; 1043(693)
g460 not 301(694) ; 1051(695)
g461 not 286(696) ; 2123(697)
g462 not 303(698) ; 1062(699)
g463 not 288(700) ; 1068(701)
g464 not 305(702) ; 1074(703)
g465 not 290(704) ; 1080(705)
g466 and 1031(630) ; 2107(706)
g467 and 1031(630) ; 2161(707)
g468 not 2154(631) ; 2158(708)
g469 and 40(29) 1387(594) 1389(610) ; 456(709)
g470 and 319(656) 36(27) 483(191) 480(292) ; 175(710)
g471 or 2036(632) 2035(519) ; 2778(711)
g472 or 2034(633) 2033(520) ; 2770(712)
g473 or 2030(637) 2029(521) ; 2754(713)
g474 or 2026(639) 2025(522) ; 2738(714)
g475 or 2038(635) 2037(523) ; 2065(715)
g476 or 2032(634) 2031(524) ; 2762(716)
g477 or 2028(638) 2027(525) ; 2746(717)
g478 or 2024(636) 2023(526) ; 2626(718)
g479 or 1751(643) 1750(527) ; 2618(719)
g480 or 1747(640) 1746(528) ; 2602(720)
g481 or 1745(641) 1744(529) ; 2594(721)
g482 or 1743(642) 1742(530) ; 2586(722)
g483 or 1739(647) 1738(531) ; 2570(723)
g484 or 1735(645) 1734(532) ; 2554(724)
g485 or 1749(644) 1748(534) ; 2610(725)
g486 or 1741(646) 1740(535) ; 2578(726)
g487 or 1737(648) 1736(536) ; 2562(727)
g488 and 1813(661) 1790(588) 1777(537) ; 1823(728)
g489 and 1536(665) 1513(593) 1500(538) ; 1546(729)
g490 or 2524(576)* 2523(653)* ; 2538(730)
g491 and 1541(577)* 1540(655)* ; 1542(731)
g492 and 1538(580)* 1537(654)* ; 1539(732)
g493 or 1234(657) 1232(659) ; 1235(733)
g494 or 2672(682)* 2665(582)* ; 2674(734)
g495 or 1227(681) 1225(660) ; 1228(735)
g496 or 2781(429)* 2778(711)* ; 2059(736)
g497 or 2773(431)* 2770(712)* ; 2055(737)
g498 or 2765(433)* 2762(716)* ; 2051(738)
g499 and 1809(662) 1786(548) 1781(574) ; 1820(739)
g500 or 2757(435)* 2754(713)* ; 2047(740)
g501 or 2749(437)* 2746(717)* ; 2043(741)
g502 or 2741(438)* 2738(714)* ; 2039(742)
g503 or 2534(663)* 2533(664)* ; 2546(743)
g504 or 2629(440)* 2626(718)* ; 1597(744)
g505 or 2621(442)* 2618(719)* ; 1593(745)
g506 or 2613(444)* 2610(725)* ; 1589(746)
g507 or 2605(446)* 2602(720)* ; 1585(747)
g508 or 2597(448)* 2594(721)* ; 1581(748)
g509 or 2589(450)* 2586(722)* ; 1577(749)
g510 and 1532(666) 1509(552) 1504(575) ; 1543(750)
g511 or 2581(452)* 2578(726)* ; 1573(751)
g512 or 2573(454)* 2570(723)* ; 1569(752)
g513 or 2565(455)* 2562(727)* ; 1565(753)
g514 or 2557(457)* 2554(724)* ; 1561(754)
g515 or 889(670) 887(597) ; 897(755)
g516 or 893(598) 891(669) ; 898(756)
g517 and 868(198) 562(672) ; 886(757)
g518 and 865(291) 562(672) ; 146(758)
g519 not 562(672) ; 2207(759)
g520 and 562(672) ; 592(760)
g521 or 2637(683)* 2634(555)* ; 1752(762)
g522 or 2645(676)* 2642(603)* ; 1761(763)
g523 or 2646(675)* 2639(605)* ; 1762(764)
g524 or 2653(678)* 2650(606)* ; 1770(765)
g525 or 2654(677)* 2647(608)* ; 1771(766)
g526 or 2661(680)* 2658(611)* ; 2663(767)
g527 or 2662(679)* 2655(613)* ; 2664(768)
g528 or 2671(658)* 2668(614)* ; 2673(769)
g529 not 2235(684) ; 2241(770)
g530 not 2110(685) ; 2114(771)
g531 not 2164(686) ; 2168(772)
g532 not 2350(687) ; 2354(773)
g533 not 2118(688) ; 2122(774)
g534 not 2262(689) ; 2266(775)
g535 not 2172(690) ; 2176(776)
g536 not 2151(691) ; 2157(777)
g537 or 2158(708)* 2151(691)* ; 2160(778)
g538 and 1043(693) ; 2342(779)
g539 and 1043(693) ; 2115(780)
g540 and 1043(693) ; 2254(781)
g541 and 1043(693) ; 2169(782)
g542 and 1051(695) ; 2422(783)
g543 and 1051(695) ; 2334(784)
g544 and 1051(695) ; 2126(785)
g545 not 2123(697) ; 2129(786)
g546 and 1062(699) ; 2134(787)
g547 and 1062(699) ; 2180(788)
g548 and 1068(701) ; 2131(789)
g549 and 1068(701) ; 2177(790)
g550 and 1074(703) ; 2144(791)
g551 and 1074(703) ; 2190(792)
g552 and 1080(705) ; 2141(793)
g553 and 1080(705) ; 2187(794)
g554 not 2107(706) ; 2113(795)
g555 not 2161(707) ; 2167(796)
g556 and 466(667) 1389(610) 40(29) ; 468(797)
g557 and 456(709) ; 995(798)
g558 not 456(709) ; 1006(799)
g559 not 456(709) ; 743(800)
g560 and 456(709) ; 749(801)
g561 not 456(709) ; 462(802)
g562 not 2778(711) ; 2782(804)
g563 not 2770(712) ; 2774(805)
g564 not 2754(713) ; 2758(806)
g565 not 2738(714) ; 2742(807)
g566 not 2762(716) ; 2766(808)
g567 not 2746(717) ; 2750(809)
g568 not 2626(718) ; 2630(810)
g569 not 2618(719) ; 2622(811)
g570 not 2602(720) ; 2606(812)
g571 not 2594(721) ; 2598(813)
g572 not 2586(722) ; 2590(814)
g573 not 2570(723) ; 2574(815)
g574 not 2554(724) ; 2558(816)
g575 not 2610(725) ; 2614(817)
g576 not 2578(726) ; 2582(818)
g577 not 2562(727) ; 2566(819)
g578 and 1821(649)* 1820(739)* ; 1822(820)
g579 and 1824(650)* 1823(728)* ; 1825(821)
g580 and 1544(651)* 1543(750)* ; 1545(822)
g581 and 1547(652)* 1546(729)* ; 1548(823)
g582 not 2538(730) ; 2542(824)
g583 or 1539(732)* 1542(731)* ; 2535(825)
g584 not 1235(733) ; 1245(826)
g585 or 2674(734)* 2673(769)* ; 2709(827)
g586 not 1228(735) ; 1243(828)
g587 or 2782(804)* 2775(341)* ; 2060(829)
g588 or 2774(805)* 2767(343)* ; 2056(830)
g589 or 2766(808)* 2759(345)* ; 2052(831)
g590 or 2758(806)* 2751(347)* ; 2048(832)
g591 or 2750(809)* 2743(350)* ; 2044(833)
g592 or 2742(807)* 2735(352)* ; 2040(834)
g593 not 2546(743) ; 2550(835)
g594 or 2630(810)* 2623(354)* ; 1598(836)
g595 or 2622(811)* 2615(356)* ; 1594(837)
g596 or 2614(817)* 2607(358)* ; 1590(838)
g597 or 2606(812)* 2599(360)* ; 1586(839)
g598 or 2598(813)* 2591(362)* ; 1582(840)
g599 or 2590(814)* 2583(364)* ; 1578(841)
g600 or 2582(818)* 2575(366)* ; 1574(842)
g601 or 2574(815)* 2567(368)* ; 1570(843)
g602 or 2566(819)* 2559(370)* ; 1566(844)
g603 or 2558(816)* 2551(372)* ; 1562(845)
g604 or 886(757) 885(596) ; 896(846)
g605 not 2207(759) ; 2213(852)
g606 not 592(760) ; 596(853)
g607 or 1753(674)* 1752(762)* ; 1754(854)
g608 and 743(800) 1701(556) ; 502(855)
g609 and 1006(799) 1701(556) ; 729(856)
g610 or 1762(764)* 1761(763)* ; 1763(857)
g611 and 743(800) 1250(604) ; 508(858)
g612 and 1006(799) 1250(604) ; 735(859)
g613 or 1771(766)* 1770(765)* ; 1772(860)
g614 or 2664(768)* 2663(767)* ; 2712(861)
g615 and 743(800) 1698(563) ; 496(862)
g616 and 1006(799) 1698(563) ; 723(863)
g617 or 2113(795)* 2110(685)* ; 569(864)
g618 or 2167(796)* 2164(686)* ; 599(865)
g619 or 2122(774)* 2115(780)* ; 579(866)
g620 or 2176(776)* 2169(782)* ; 609(867)
g621 not 2342(779) ; 2346(868)
g622 not 2115(780) ; 2121(869)
g623 not 2254(781) ; 2258(870)
g624 not 2169(782) ; 2175(871)
g625 not 2422(783) ; 2426(872)
g626 not 2334(784) ; 2338(873)
g627 or 2129(786)* 2126(785)* ; 587(874)
g628 not 2126(785) ; 2130(875)
g629 and 749(801) 286(696) ; 765(876)
g630 and 995(798) 286(696) ; 1014(877)
g631 and 749(801) 303(698) ; 769(878)
g632 and 995(798) 303(698) ; 1018(879)
g633 not 2134(787) ; 2138(880)
g634 not 2180(788) ; 2184(881)
g635 not 2131(789) ; 2137(882)
g636 not 2177(790) ; 2183(883)
g637 not 2144(791) ; 2148(884)
g638 not 2190(792) ; 2194(885)
g639 and 743(800) 290(704) ; 490(886)
g640 and 1006(799) 290(704) ; 717(887)
g641 not 2141(793) ; 2147(888)
g642 not 2187(794) ; 2193(889)
g643 or 2114(771)* 2107(706)* ; 570(890)
g644 or 2168(772)* 2161(707)* ; 600(891)
g645 or 2157(777)* 2154(631)* ; 2159(892)
g646 and 468(797) ; 1257(893)
g647 and 468(797) ; 1258(894)
g648 not 995(798) ; 999(895)
g649 not 749(801) ; 753(896)
g650 and 462(802) ; 475(897)
g651 and 462(802) ; 1337(898)
g652 or 1822(820)* 1825(821)* ; 2727(899)
g653 or 1545(822)* 1548(823)* ; 2543(900)
g654 or 2542(824)* 2535(825)* ; 1550(901)
g655 not 2535(825) ; 2541(902)
g656 and 1245(826) 1235(733) ; 1094(903)
g657 not 2709(827) ; 2715(904)
g658 and 1243(828) 1228(735) ; 1096(905)
g659 or 2060(829)* 2059(736)* ; 2061(906)
g660 or 2056(830)* 2055(737)* ; 2057(907)
g661 or 2052(831)* 2051(738)* ; 2053(908)
g662 or 2048(832)* 2047(740)* ; 2049(909)
g663 or 2044(833)* 2043(741)* ; 2045(910)
g664 or 2040(834)* 2039(742)* ; 2041(911)
g665 or 1598(836)* 1597(744)* ; 1599(912)
g666 or 1594(837)* 1593(745)* ; 1595(913)
g667 or 1590(838)* 1589(746)* ; 1591(914)
g668 or 1586(839)* 1585(747)* ; 1587(915)
g669 or 1582(840)* 1581(748)* ; 1583(916)
g670 or 1578(841)* 1577(749)* ; 1579(917)
g671 or 1574(842)* 1573(751)* ; 1575(918)
g672 or 1570(843)* 1569(752)* ; 1571(919)
g673 or 1566(844)* 1565(753)* ; 1567(920)
g674 or 1562(845)* 1561(754)* ; 1563(921)
g675 not 1754(854) ; 1758(924)
g676 not 1763(857) ; 1767(925)
g677 and 1772(860) ; 1802(926)
g678 and 1772(860) ; 1798(927)
g679 not 2712(861) ; 2716(928)
g680 or 570(890)* 569(864)* ; 571(929)
g681 or 600(891)* 599(865)* ; 601(930)
g682 or 2121(869)* 2118(688)* ; 578(931)
g683 or 2175(871)* 2172(690)* ; 608(932)
g684 or 2160(778)* 2159(892)* ; 2210(933)
g685 and 753(896) 286(696) ; 763(934)
g686 and 999(895) 286(696) ; 1012(935)
g687 or 2130(875)* 2123(697)* ; 588(936)
g688 and 753(896) 303(698) ; 767(937)
g689 and 999(895) 303(698) ; 1016(938)
g690 or 2137(882)* 2134(787)* ; 2139(939)
g691 or 2183(883)* 2180(788)* ; 2185(940)
g692 and 753(896) 288(700) ; 531(941)
g693 and 999(895) 288(700) ; 705(942)
g694 or 2138(880)* 2131(789)* ; 2140(943)
g695 or 2184(881)* 2177(790)* ; 2186(944)
g696 and 753(896) 305(702) ; 537(945)
g697 and 999(895) 305(702) ; 711(946)
g698 or 2147(888)* 2144(791)* ; 2149(947)
g699 or 2193(889)* 2190(792)* ; 2195(948)
g700 or 2148(884)* 2141(793)* ; 2150(949)
g701 or 2194(885)* 2187(794)* ; 2196(950)
g702 and 1257(893) ; 742(951)
g703 and 1257(893) ; 1005(952)
g704 and 1258(894) ; 1845(953)
g705 and 1258(894) ; 1907(954)
g706 and 475(897) ; 1836(955)
g707 and 475(897) ; 1850(956)
g708 and 475(897) ; 1355(957)
g709 and 1337(898) ; 1898(958)
g710 and 1337(898) ; 1912(959)
g711 and 1337(898) ; 1601(960)
g712 not 2727(899) ; 2733(961)
g713 not 2543(900) ; 2549(962)
g714 or 2541(902)* 2538(730)* ; 1549(963)
g715 or 1245(826) 1094(903) ; 154(964)
g716 or 2716(928)* 2709(827)* ; 2718(965)
g717 or 2734(584)* 2727(899)* ; 1829(966)
g718 or 1243(828) 1096(905) ; 155(967)
g719 not 2061(906) ; 2062(968)
g720 not 2057(907) ; 2058(969)
g721 not 2053(908) ; 2054(970)
g722 not 2049(909) ; 2050(971)
g723 and 1850(956) 2070(260) ; 1876(972)
g724 and 1912(959) 2070(260) ; 1938(973)
g725 not 2045(910) ; 2046(974)
g726 and 1850(956) 1999(265) ; 1874(975)
g727 and 1912(959) 1999(265) ; 1936(976)
g728 not 2041(911) ; 2042(977)
g729 or 2550(835)* 2543(900)* ; 1552(978)
g730 and 1850(956) 1994(267) ; 1872(979)
g731 and 1912(959) 1994(267) ; 1934(980)
g732 not 1599(912) ; 1600(981)
g733 and 1850(956) 1989(269) ; 1870(982)
g734 and 1912(959) 1989(269) ; 1932(983)
g735 not 1595(913) ; 1596(984)
g736 and 1836(955) 1984(271) ; 1868(985)
g737 and 1898(958) 1984(271) ; 1930(986)
g738 not 1591(914) ; 1592(987)
g739 and 1836(955) 1979(273) ; 1866(988)
g740 and 1898(958) 1979(273) ; 1928(989)
g741 not 1587(915) ; 1588(990)
g742 and 1836(955) 1974(275) ; 1863(991)
g743 and 1898(958) 1974(275) ; 1925(992)
g744 not 1583(916) ; 1584(993)
g745 and 1836(955) 1969(277) ; 1858(994)
g746 and 1898(958) 1969(277) ; 1920(995)
g747 not 1579(917) ; 1580(996)
g748 and 1355(957) 1964(279) ; 1377(997)
g749 and 1601(960) 1964(279) ; 1623(998)
g750 not 1575(918) ; 1576(999)
g751 and 1355(957) 1959(281) ; 1373(1000)
g752 and 1601(960) 1959(281) ; 1619(1001)
g753 not 1571(919) ; 1572(1002)
g754 and 1601(960) 1351(284) ; 1615(1003)
g755 and 1355(957) 1351(284) ; 1369(1004)
g756 not 1567(920) ; 1568(1005)
g757 and 1355(957) 1344(286) ; 676(1006)
g758 and 1601(960) 1344(286) ; 1108(1007)
g759 not 1563(921) ; 1564(1008)
g760 or 2213(852)* 2210(933)* ; 2215(1009)
g761 and 1798(927) 1754(854) 1763(857) ; 1815(1010)
g762 and 1802(926) 1758(924) 1767(925) ; 1818(1011)
g763 and 742(951) 502(855) ; 504(1012)
g764 and 1005(952) 729(856) ; 731(1013)
g765 and 742(951) 508(858) ; 510(1014)
g766 and 1005(952) 735(859) ; 737(1015)
g767 not 1802(926) ; 1805(1016)
g768 not 1798(927) ; 1801(1017)
g769 or 2715(904)* 2712(861)* ; 2717(1018)
g770 and 742(951) 496(862) ; 498(1019)
g771 and 1005(952) 723(863) ; 725(1020)
g772 not 571(929) ; 575(1021)
g773 not 601(930) ; 605(1022)
g774 or 579(866)* 578(931)* ; 580(1023)
g775 or 609(867)* 608(932)* ; 610(1024)
g776 not 2210(933) ; 2214(1025)
g777 or 588(936)* 587(874)* ; 589(1026)
g778 or 765(876) 763(934) ; 519(1027)
g779 or 1014(877) 1012(935) ; 693(1028)
g780 or 769(878) 767(937) ; 525(1029)
g781 or 1018(879) 1016(938) ; 699(1030)
g782 or 2140(943)* 2139(939)* ; 2200(1031)
g783 or 2186(944)* 2185(940)* ; 2220(1032)
g784 or 2150(949)* 2149(947)* ; 2197(1033)
g785 or 2196(950)* 2195(948)* ; 2217(1034)
g786 and 742(951) 490(886) ; 492(1035)
g787 and 1005(952) 717(887) ; 719(1036)
g788 not 1836(955) ; 1842(1037)
g789 not 1355(957) ; 1361(1038)
g790 not 1898(958) ; 1904(1039)
g791 not 1601(960) ; 1607(1040)
g792 and 748(411) 531(941) ; 533(1041)
g793 and 748(411) 537(945) ; 539(1042)
g794 and 994(412) 705(942) ; 707(1043)
g795 and 994(412) 711(946) ; 713(1044)
g796 or 1550(901)* 1549(963)* ; 1091(1045)
g797 or 2718(965)* 2717(1018)* ; 2722(1047)
g798 or 2733(961)* 2730(546)* ; 1828(1048)
g799 and 1842(1037) 2094(251) ; 1861(1049)
g800 and 1904(1039) 2094(251) ; 1923(1050)
g801 and 1842(1037) 2088(253) ; 1856(1051)
g802 and 1904(1039) 2088(253) ; 1918(1052)
g803 and 2042(977) 2046(974) 2050(971) 2054(970) 2058(969) ; 1558(1053)
g804 and 1361(1038) 2082(255) ; 1375(1054)
g805 and 1607(1040) 2082(255) ; 1621(1055)
g806 and 1361(1038) 2076(257) ; 1371(1056)
g807 and 1607(1040) 2076(257) ; 1617(1057)
g808 and 1361(1038) 2070(260) ; 1368(1058)
g809 and 1607(1040) 2070(260) ; 1614(1059)
g810 and 1361(1038) 1999(265) ; 675(1060)
g811 and 1607(1040) 1999(265) ; 1107(1061)
g812 or 2549(962)* 2546(743)* ; 1551(1062)
g813 and 1584(993) 1588(990) 1592(987) 1596(984) 1600(981) ; 1554(1063)
g814 and 1564(1008) 1568(1005) 1572(1002) 1576(999) 1580(996) ; 1555(1064)
g815 or 2214(1025)* 2207(759)* ; 2216(1065)
g816 and 1805(1016) 1767(925) 1754(854) ; 1817(1066)
g817 not 504(1012) ; 505(1067)
g818 not 731(1013) ; 732(1068)
g819 and 1801(1017) 1763(857) 1758(924) ; 1814(1069)
g820 not 510(1014) ; 511(1070)
g821 not 737(1015) ; 738(1071)
g822 not 498(1019) ; 499(1072)
g823 not 725(1020) ; 726(1073)
g824 not 580(1023) ; 584(1074)
g825 and 610(1024) ; 621(1075)
g826 and 610(1024) ; 625(1076)
g827 and 589(1026) ; 617(1077)
g828 and 589(1026) ; 613(1078)
g829 not 2200(1031) ; 2204(1079)
g830 not 2220(1032) ; 2224(1080)
g831 not 2197(1033) ; 2203(1081)
g832 not 2217(1034) ; 2223(1082)
g833 not 492(1035) ; 493(1083)
g834 not 719(1036) ; 720(1084)
g835 and 1845(953) 1874(975) ; 1889(1085)
g836 and 1845(953) 1872(979) ; 1887(1086)
g837 and 1845(953) 1870(982) ; 1885(1087)
g838 and 1845(953) 1876(972) ; 1891(1088)
g839 and 1907(954) 1936(976) ; 1951(1089)
g840 and 1907(954) 1934(980) ; 1949(1090)
g841 and 1907(954) 1932(983) ; 1947(1091)
g842 and 1907(954) 1938(973) ; 1953(1092)
g843 and 2062(968) 2065(715) ; 1557(1093)
g844 and 1831(409) 1868(985) ; 1883(1094)
g845 and 1831(409) 1866(988) ; 1881(1095)
g846 and 1893(410) 1930(986) ; 1945(1096)
g847 and 1893(410) 1928(989) ; 1943(1097)
g848 and 748(411) 519(1027) ; 521(1098)
g849 and 748(411) 525(1029) ; 527(1099)
g850 not 533(1041) ; 534(1100)
g851 not 539(1042) ; 540(1101)
g852 and 994(412) 693(1028) ; 695(1102)
g853 and 994(412) 699(1030) ; 701(1103)
g854 not 707(1043) ; 708(1104)
g855 not 713(1044) ; 714(1105)
g856 not 1091(1045) ; 1092(1106)
g857 not 2722(1047) ; 2726(1107)
g858 or 1829(966)* 1828(1048)* ; 1830(1108)
g859 and 1558(1053) 1557(1093) ; 1559(1109)
g860 or 1552(978)* 1551(1062)* ; 1553(1110)
g861 and 1555(1064) 1554(1063) ; 1556(1111)
g862 or 1863(991) 1861(1049) ; 1864(1112)
g863 or 1925(992) 1923(1050) ; 1926(1113)
g864 or 1858(994) 1856(1051) ; 1859(1114)
g865 or 1920(995) 1918(1052) ; 1921(1115)
g866 or 1377(997) 1375(1054) ; 1382(1116)
g867 or 1623(998) 1621(1055) ; 1628(1117)
g868 or 1373(1000) 1371(1056) ; 1380(1118)
g869 or 1619(1001) 1617(1057) ; 1626(1119)
g870 or 1615(1003) 1614(1059) ; 1624(1120)
g871 or 1369(1004) 1368(1058) ; 1378(1121)
g872 or 676(1006) 675(1060) ; 677(1122)
g873 or 1108(1007) 1107(1061) ; 1109(1123)
g874 or 2216(1065)* 2215(1009)* ; 2238(1124)
g875 and 621(1075) 592(760) 601(930) ; 636(1125)
g876 and 625(1076) 596(853) 605(1022) ; 639(1126)
g877 and 1815(1010)* 1814(1069)* ; 1816(1127)
g878 and 1818(1011)* 1817(1066)* ; 1819(1128)
g879 and 505(1067) 1889(1085) ; 915(1129)
g880 and 505(1067) ; 2278(1130)
g881 and 732(1068) 1951(1089) ; 1133(1131)
g882 and 732(1068) ; 2366(1132)
g883 and 511(1070) 1891(1088) ; 907(1133)
g884 and 511(1070) ; 2270(1134)
g885 and 738(1071) 1953(1092) ; 1125(1135)
g886 and 738(1071) ; 2358(1136)
g887 and 499(1072) 1887(1086) ; 922(1137)
g888 and 499(1072) ; 2286(1138)
g889 and 726(1073) 1949(1090) ; 1140(1139)
g890 and 726(1073) ; 2374(1140)
g891 and 613(1078) 571(929) 580(1023) ; 630(1141)
g892 and 617(1077) 575(1021) 584(1074) ; 633(1142)
g893 not 621(1075) ; 624(1143)
g894 not 625(1076) ; 628(1144)
g895 not 617(1077) ; 620(1145)
g896 not 613(1078) ; 616(1146)
g897 or 2203(1081)* 2200(1031)* ; 2205(1147)
g898 or 2223(1082)* 2220(1032)* ; 2225(1148)
g899 or 2204(1079)* 2197(1033)* ; 2206(1149)
g900 or 2224(1080)* 2217(1034)* ; 2226(1150)
g901 and 1885(1087) 493(1083) ; 924(1151)
g902 and 493(1083) ; 2294(1152)
g903 and 1947(1091) 720(1084) ; 1142(1153)
g904 and 720(1084) ; 2382(1154)
g905 and 1889(1085) ; 2275(1155)
g906 and 1887(1086) ; 2283(1156)
g907 and 1885(1087) ; 2291(1157)
g908 and 1891(1088) ; 2267(1158)
g909 and 1951(1089) ; 2363(1159)
g910 and 1949(1090) ; 2371(1160)
g911 and 1947(1091) ; 2379(1161)
g912 and 1953(1092) ; 2355(1162)
g913 and 540(1101) 1883(1094) ; 937(1163)
g914 and 1883(1094) ; 2299(1164)
g915 and 534(1100) 1881(1095) ; 946(1165)
g916 and 1881(1095) ; 2307(1166)
g917 and 714(1105) 1945(1096) ; 1155(1167)
g918 and 1945(1096) ; 2387(1168)
g919 and 708(1104) 1943(1097) ; 1164(1169)
g920 and 1943(1097) ; 2395(1170)
g921 not 521(1098) ; 522(1171)
g922 not 527(1099) ; 528(1172)
g923 and 534(1100) ; 2310(1173)
g924 and 540(1101) ; 2302(1174)
g925 not 695(1102) ; 696(1175)
g926 not 701(1103) ; 702(1176)
g927 and 708(1104) ; 2398(1177)
g928 and 714(1105) ; 2390(1178)
g929 and 1382(1116) ; 2331(1181)
g930 and 1628(1117) ; 2419(1182)
g931 and 1380(1118) ; 2251(1183)
g932 and 1626(1119) ; 2339(1184)
g933 and 1624(1120) ; 2347(1185)
g934 and 1378(1121) ; 2259(1186)
g935 not 2238(1124) ; 2242(1187)
g936 and 628(1144) 605(1022) 592(760) ; 638(1188)
g937 and 624(1143) 601(930) 596(853) ; 635(1189)
g938 or 1816(1127)* 1819(1128)* ; 2719(1190)
g939 not 2278(1130) ; 2282(1191)
g940 not 2366(1132) ; 2370(1192)
g941 not 2270(1134) ; 2274(1193)
g942 not 2358(1136) ; 2362(1194)
g943 not 2286(1138) ; 2290(1195)
g944 not 2374(1140) ; 2378(1196)
g945 or 2241(770)* 2238(1124)* ; 645(1197)
g946 and 620(1145) 584(1074) 571(929) ; 632(1198)
g947 and 616(1146) 580(1023) 575(1021) ; 629(1199)
g948 and 1035(618) 1378(1121) ; 674(1200)
g949 and 1035(618) 1624(1120) ; 1106(1201)
g950 and 1043(693) 1380(1118) ; 671(1202)
g951 and 1043(693) 1626(1119) ; 1104(1203)
g952 and 1051(695) 1382(1116) ; 967(1204)
g953 and 1051(695) 1628(1117) ; 1184(1205)
g954 or 2206(1149)* 2205(1147)* ; 2230(1206)
g955 or 2226(1150)* 2225(1148)* ; 2246(1207)
g956 not 2294(1152) ; 2298(1208)
g957 not 2382(1154) ; 2386(1209)
g958 and 1031(630) 677(1122) ; 679(1210)
g959 and 1031(630) 1109(1123) ; 1110(1211)
g960 not 2275(1155) ; 2281(1212)
g961 not 2283(1156) ; 2289(1213)
g962 not 2291(1157) ; 2297(1214)
g963 not 2267(1158) ; 2273(1215)
g964 not 2363(1159) ; 2369(1216)
g965 not 2371(1160) ; 2377(1217)
g966 not 2379(1161) ; 2385(1218)
g967 not 2355(1162) ; 2361(1219)
g968 and 14(9) 1092(1106) ; 401(1276)
g969 and 894(533) 1559(1109) 1556(1111) ; 311(1278)
g970 not 2299(1164) ; 2305(1222)
g971 not 2307(1166) ; 2313(1223)
g972 and 1831(409) 1864(1112) ; 1879(1224)
g973 and 1831(409) 1859(1114) ; 1877(1225)
g974 not 2387(1168) ; 2393(1226)
g975 not 2395(1170) ; 2401(1227)
g976 and 1893(410) 1926(1113) ; 1941(1228)
g977 and 1893(410) 1921(1115) ; 1939(1229)
g978 and 522(1171) ; 2326(1230)
g979 and 528(1172) ; 2318(1231)
g980 not 2310(1173) ; 2314(1232)
g981 not 2302(1174) ; 2306(1233)
g982 and 696(1175) ; 2414(1234)
g983 and 702(1176) ; 2406(1235)
g984 not 2398(1177) ; 2402(1236)
g985 not 2390(1178) ; 2394(1237)
g986 or 2726(1107)* 2719(1190)* ; 1827(1238)
g987 not 2331(1181) ; 2337(1239)
g988 not 2419(1182) ; 2425(1240)
g989 not 2251(1183) ; 2257(1241)
g990 not 2339(1184) ; 2345(1242)
g991 not 2347(1185) ; 2353(1243)
g992 not 2259(1186) ; 2265(1244)
g993 and 636(1125)* 635(1189)* ; 637(1245)
g994 and 639(1126)* 638(1188)* ; 640(1246)
g995 not 2719(1190) ; 2725(1247)
g996 or 2281(1212)* 2278(1130)* ; 908(1248)
g997 or 2369(1216)* 2366(1132)* ; 1126(1249)
g998 or 2273(1215)* 2270(1134)* ; 899(1250)
g999 or 2361(1219)* 2358(1136)* ; 1117(1251)
g1000 or 2289(1213)* 2286(1138)* ; 916(1252)
g1001 or 2377(1217)* 2374(1140)* ; 1134(1253)
g1002 or 2242(1187)* 2235(684)* ; 646(1254)
g1003 and 630(1141)* 629(1199)* ; 631(1255)
g1004 and 633(1142)* 632(1198)* ; 634(1256)
g1005 or 2354(773)* 2347(1185)* ; 1115(1257)
g1006 or 2266(775)* 2259(1186)* ; 684(1258)
g1007 or 2346(868)* 2339(1184)* ; 1099(1259)
g1008 or 2258(870)* 2251(1183)* ; 665(1260)
g1009 or 2426(872)* 2419(1182)* ; 1181(1261)
g1010 or 2338(873)* 2331(1181)* ; 963(1262)
g1011 not 2230(1206) ; 2234(1263)
g1012 not 2246(1207) ; 2250(1264)
g1013 or 2297(1214)* 2294(1152)* ; 925(1265)
g1014 or 2385(1218)* 2382(1154)* ; 1143(1266)
g1015 or 2282(1191)* 2275(1155)* ; 909(1267)
g1016 or 2290(1195)* 2283(1156)* ; 917(1268)
g1017 or 2298(1208)* 2291(1157)* ; 926(1269)
g1018 or 2274(1193)* 2267(1158)* ; 900(1270)
g1019 or 2370(1192)* 2363(1159)* ; 1127(1271)
g1020 or 2378(1196)* 2371(1160)* ; 1135(1272)
g1021 or 2386(1209)* 2379(1161)* ; 1144(1273)
g1022 or 2362(1194)* 2355(1162)* ; 1118(1274)
g1023 not 401(1276) ; 1087(1275)
g1024 or 2306(1233)* 2299(1164)* ; 929(1279)
g1025 or 2314(1232)* 2307(1166)* ; 939(1280)
g1026 and 1879(1224) ; 2315(1281)
g1027 and 1877(1225) ; 2323(1282)
g1028 or 2394(1237)* 2387(1168)* ; 1147(1283)
g1029 or 2402(1236)* 2395(1170)* ; 1157(1284)
g1030 and 1941(1228) ; 2403(1285)
g1031 and 1939(1229) ; 2411(1286)
g1032 not 2326(1230) ; 2330(1287)
g1033 and 522(1171) 1877(1225) ; 961(1288)
g1034 and 528(1172) 1879(1224) ; 954(1289)
g1035 not 2318(1231) ; 2322(1290)
g1036 or 2313(1223)* 2310(1173)* ; 938(1291)
g1037 or 2305(1222)* 2302(1174)* ; 928(1292)
g1038 not 2414(1234) ; 2418(1293)
g1039 and 696(1175) 1939(1229) ; 1179(1294)
g1040 and 702(1176) 1941(1228) ; 1172(1295)
g1041 not 2406(1235) ; 2410(1296)
g1042 or 2401(1227)* 2398(1177)* ; 1156(1297)
g1043 or 2393(1226)* 2390(1178)* ; 1146(1298)
g1044 or 2725(1247)* 2722(1047)* ; 1826(1299)
g1045 or 637(1245)* 640(1246)* ; 2243(1300)
g1046 or 909(1267)* 908(1248)* ; 910(1301)
g1047 or 1127(1271)* 1126(1249)* ; 1128(1302)
g1048 or 900(1270)* 899(1250)* ; 901(1303)
g1049 or 1118(1274)* 1117(1251)* ; 1119(1304)
g1050 or 917(1268)* 916(1252)* ; 918(1305)
g1051 or 1135(1272)* 1134(1253)* ; 1136(1306)
g1052 or 646(1254)* 645(1197)* ; 647(1307)
g1053 or 631(1255)* 634(1256)* ; 2227(1308)
g1054 or 2353(1243)* 2350(687)* ; 1114(1309)
g1055 or 2265(1244)* 2262(689)* ; 683(1310)
g1056 or 2345(1242)* 2342(779)* ; 1098(1311)
g1057 or 2257(1241)* 2254(781)* ; 664(1312)
g1058 or 2425(1240)* 2422(783)* ; 1180(1313)
g1059 or 2337(1239)* 2334(784)* ; 962(1314)
g1060 or 926(1269)* 925(1265)* ; 927(1315)
g1061 or 1144(1273)* 1143(1266)* ; 1145(1316)
g1062 or 929(1279)* 928(1292)* ; 930(1317)
g1063 or 939(1280)* 938(1291)* ; 940(1318)
g1064 or 2322(1290)* 2315(1281)* ; 948(1319)
g1065 not 2315(1281) ; 2321(1320)
g1066 or 2330(1287)* 2323(1282)* ; 956(1321)
g1067 not 2323(1282) ; 2329(1322)
g1068 or 1147(1283)* 1146(1298)* ; 1148(1323)
g1069 or 1157(1284)* 1156(1297)* ; 1158(1324)
g1070 or 2410(1296)* 2403(1285)* ; 1166(1325)
g1071 not 2403(1285) ; 2409(1326)
g1072 or 2418(1293)* 2411(1286)* ; 1174(1327)
g1073 not 2411(1286) ; 2417(1328)
g1074 or 1827(1238)* 1826(1299)* ; 686(1329)
g1075 and 865(291) 647(1307) ; 143(1330)
g1076 not 2243(1300) ; 2249(1331)
g1077 and 915(1129) 901(1303) ; 970(1332)
g1078 and 901(1303) 918(1305) 927(1315) 910(1301) ; 968(1333)
g1079 and 1133(1131) 1119(1304) ; 1187(1334)
g1080 and 1119(1304) 1136(1306) 1145(1316) 1128(1302) ; 1185(1335)
g1081 and 922(1137) 901(1303) 910(1301) ; 971(1336)
g1082 and 1140(1139) 1119(1304) 1128(1302) ; 1188(1337)
g1083 not 2227(1308) ; 2233(1338)
g1084 or 1115(1257)* 1114(1309)* ; 1112(1339)
g1085 or 684(1258)* 683(1310)* ; 681(1340)
g1086 or 1099(1259)* 1098(1311)* ; 1100(1341)
g1087 or 665(1260)* 664(1312)* ; 666(1342)
g1088 or 1181(1261)* 1180(1313)* ; 1182(1343)
g1089 or 963(1262)* 962(1314)* ; 964(1344)
g1090 or 2234(1263)* 2227(1308)* ; 642(1345)
g1091 or 2250(1264)* 2243(1300)* ; 649(1346)
g1092 and 910(1301) 924(1151) 901(1303) 918(1305) ; 972(1347)
g1093 and 1128(1302) 1142(1153) 1119(1304) 1136(1306) ; 1189(1348)
g1094 and 946(1165) 930(1317) ; 978(1349)
g1095 and 1164(1169) 1148(1323) ; 1195(1350)
g1096 or 2329(1322)* 2326(1230)* ; 955(1351)
g1097 and 954(1289) 930(1317) 940(1318) ; 979(1352)
g1098 or 2321(1320)* 2318(1231)* ; 947(1353)
g1099 or 2417(1328)* 2414(1234)* ; 1173(1354)
g1100 and 1172(1295) 1148(1323) 1158(1324) ; 1196(1355)
g1101 or 2409(1326)* 2406(1235)* ; 1165(1356)
g1102 not 686(1329) ; 687(1357)
g1103 not 968(1333) ; 969(1359)
g1104 not 1185(1335) ; 1186(1360)
g1105 or 972(1347) 971(1336) 970(1332) 907(1133) ; 973(1361)
g1106 or 1189(1348) 1188(1337) 1187(1334) 1125(1135) ; 1190(1362)
g1107 and 674(1200) 666(1342) ; 680(1363)
g1108 and 1106(1201) 1100(1341) ; 1111(1364)
g1109 or 2233(1338)* 2230(1206)* ; 641(1365)
g1110 or 2249(1331)* 2246(1207)* ; 648(1366)
g1111 and 679(1210) 666(1342) 681(1340) ; 682(1367)
g1112 and 1110(1211) 1100(1341) 1112(1339) ; 1113(1368)
g1113 or 948(1319)* 947(1353)* ; 949(1369)
g1114 or 956(1321)* 955(1351)* ; 957(1370)
g1115 or 1166(1325)* 1165(1356)* ; 1167(1371)
g1116 or 1174(1327)* 1173(1354)* ; 1175(1372)
g1117 not 973(1361) ; 976(1373)
g1118 not 1190(1362) ; 1193(1374)
g1119 or 682(1367) 680(1363) 671(1202) ; 685(1375)
g1120 or 1113(1368) 1111(1364) 1104(1203) ; 1116(1376)
g1121 and 940(1318) 967(1204) 930(1317) 949(1369) 957(1370) ; 981(1377)
g1122 and 1158(1324) 1184(1205) 1148(1323) 1167(1371) 1175(1372) ; 1198(1378)
g1123 or 642(1345)* 641(1365)* ; 643(1379)
g1124 or 649(1346)* 648(1366)* ; 650(1380)
g1125 and 487(403) 687(1357) ; 395(1392)
g1126 and 957(1370) 930(1317) 949(1369) 964(1344) 940(1318) ; 977(1382)
g1127 and 1175(1372) 1148(1323) 1167(1371) 1182(1343) 1158(1324) ; 1194(1383)
g1128 and 940(1318) 961(1288) 930(1317) 949(1369) ; 980(1384)
g1129 and 1158(1324) 1179(1294) 1148(1323) 1167(1371) ; 1197(1385)
g1130 and 868(198) 650(1380) ; 884(1386)
g1131 or 969(1359)* 976(1373)* ; 988(1387)
g1132 or 1186(1360)* 1193(1374)* ; 1205(1388)
g1133 and 685(1375) 977(1382) ; 983(1389)
g1134 and 1116(1376) 1194(1383) ; 1200(1390)
g1135 not 643(1379) ; 644(1391)
g1136 not 395(1392) ; 690(1393)
g1137 or 981(1377) 980(1384) 979(1352) 978(1349) 937(1163) ; 982(1394)
g1138 or 1198(1378) 1197(1385) 1196(1355) 1195(1350) 1155(1167) ; 1199(1395)
g1139 or 884(1386) 883(668) ; 895(1396)
g1140 or 983(1389) 982(1394) ; 984(1397)
g1141 or 1200(1390) 1199(1395) ; 1201(1398)
g1142 and 487(403) 644(1391) ; 397(1406)
g1143 and 984(1397) 988(1387) ; 990(1402)
g1144 and 1201(1398) 1205(1388) ; 1207(1403)
g1145 not 984(1397) ; 987(1404)
g1146 not 1201(1398) ; 1204(1405)
g1147 not 397(1406) ; 1027(1407)
g1148 and 1830(1108) 1027(1407) 690(1393) ; 1085(1408)
g1149 and 987(1404) 973(1361) ; 989(1409)
g1150 and 1204(1405) 1190(1362) ; 1206(1410)
g1151 or 990(1402) 989(1409) ; 991(1411)
g1152 or 1207(1403) 1206(1410) ; 329(1414)
g1153 or 991(1411)* 329(1414)* ; 1221(1413)
g1154 and 991(1411) 1221(1413) ; 1239(1415)
g1155 and 1221(1413) 329(1414) ; 1238(1416)
g1156 or 1239(1415) 1238(1416) ; 1240(1417)
g1157 not 1240(1417) ; 1247(1418)
g1158 and 1247(1418) 1240(1417) ; 471(1419)
g1159 or 1247(1418) 471(1419) ; 473(1420)
g1160 and 473(1420) 1087(1275) 1553(1110) ; 1088(1421)
g1161 and 319(656) 1088(1421) 1085(1408) ; 308(1425)
g1162 and IN-169(114) ; 169(114)
g1163 and IN-174(115) ; 174(115)
g1164 and IN-177(116) ; 177(116)
g1165 and IN-178(117) ; 178(117)
g1166 and IN-179(118) ; 179(118)
g1167 and IN-180(119) ; 180(119)
g1168 and IN-181(120) ; 181(120)
g1169 and IN-182(121) ; 182(121)
g1170 and IN-183(122) ; 183(122)
g1171 and IN-184(123) ; 184(123)
g1172 and IN-185(124) ; 185(124)
g1173 and IN-186(125) ; 186(125)
g1174 and IN-189(126) ; 189(126)
g1175 and IN-190(127) ; 190(127)
g1176 and IN-191(128) ; 191(128)
g1177 and IN-192(129) ; 192(129)
g1178 and IN-193(130) ; 193(130)
g1179 and IN-194(131) ; 194(131)
g1180 and IN-195(132) ; 195(132)
g1181 and IN-196(133) ; 196(133)
g1182 and IN-197(134) ; 197(134)
g1183 and IN-198(135) ; 198(135)
g1184 and IN-199(136) ; 199(136)
g1185 and IN-200(137) ; 200(137)
g1186 and IN-201(138) ; 201(138)
g1187 and IN-202(139) ; 202(139)
g1188 and IN-203(140) ; 203(140)
g1189 and IN-204(141) ; 204(141)
g1190 and IN-205(142) ; 205(142)
g1191 and IN-206(143) ; 206(143)
g1192 and IN-207(144) ; 207(144)
g1193 and IN-208(145) ; 208(145)
g1194 and IN-209(146) ; 209(146)
g1195 and IN-210(147) ; 210(147)
g1196 and IN-211(148) ; 211(148)
g1197 and IN-212(149) ; 212(149)
g1198 and IN-213(150) ; 213(150)
g1199 and IN-214(151) ; 214(151)
g1200 and IN-215(152) ; 215(152)
g1201 and IN-239(153) ; 239(153)
g1202 and IN-240(154) ; 240(154)
g1203 and IN-241(155) ; 241(155)
g1204 and IN-242(156) ; 242(156)
g1205 and IN-243(157) ; 243(157)
g1206 and IN-244(158) ; 244(158)
g1207 and IN-245(159) ; 245(159)
g1208 and IN-246(160) ; 246(160)
g1209 and IN-247(161) ; 247(161)
g1210 and IN-248(162) ; 248(162)
g1211 and IN-249(163) ; 249(163)
g1212 and IN-250(164) ; 250(164)
g1213 and IN-251(165) ; 251(165)
g1214 and IN-252(166) ; 252(166)
g1215 and IN-253(167) ; 253(167)
g1216 and IN-254(168) ; 254(168)
g1217 and IN-255(169) ; 255(169)
g1218 and IN-256(170) ; 256(170)
g1219 and IN-257(171) ; 257(171)
g1220 and IN-262(172) ; 262(172)
g1221 and IN-263(173) ; 263(173)
g1222 and IN-264(174) ; 264(174)
g1223 and IN-265(175) ; 265(175)
g1224 and IN-266(176) ; 266(176)
g1225 and IN-267(177) ; 267(177)
g1226 and IN-268(178) ; 268(178)
g1227 and IN-269(179) ; 269(179)
g1228 and IN-270(180) ; 270(180)
g1229 and IN-271(181) ; 271(181)
g1230 and IN-272(182) ; 272(182)
g1231 and IN-273(183) ; 273(183)
g1232 and IN-274(184) ; 274(184)
g1233 and IN-275(185) ; 275(185)
g1234 and IN-276(186) ; 276(186)
g1235 and IN-277(187) ; 277(187)
g1236 and IN-278(188) ; 278(188)
g1237 and IN-279(189) ; 279(189)
g1238 and 452(190) ; 350(301)
g1239 and 452(190) ; 335(299)
g1240 and 452(190) ; 409(298)
g1241 and 1083(199) ; 369(289)
g1242 and 1083(199) ; 367(288)
g1243 and 2066(212) ; 411(264)
g1244 and 2066(212) ; 337(263)
g1245 and 2066(212) ; 384(262)
g1246 and 897(755) ; 284(847)
g1247 and 897(755) ; 321(848)
g1248 and 898(756) ; 297(849)
g1249 and 898(756) ; 280(850)
g1250 and 896(846) ; 282(922)
g1251 and 896(846) ; 323(923)
g1252 and 895(1396) ; 295(1400)
g1253 and 895(1396) ; 331(1401)
g1254 not 567(194) ; 567(194)*
g1255 not 1955(320) ; 1955(320)*
g1256 not 154(964) ; 154(964)*
g1257 not 155(967) ; 155(967)*
g1258 not 2675(261) ; 2675(261)*
g1259 not 2682(233) ; 2682(233)*
g1260 not 2471(282) ; 2471(282)*
g1261 not 2478(234) ; 2478(234)*
g1262 not 2454(230) ; 2454(230)*
g1263 not 2457(236) ; 2457(236)*
g1264 not 2451(229) ; 2451(229)*
g1265 not 2458(235) ; 2458(235)*
g1266 not 2446(228) ; 2446(228)*
g1267 not 2449(238) ; 2449(238)*
g1268 not 2443(227) ; 2443(227)*
g1269 not 2450(237) ; 2450(237)*
g1270 not 2438(226) ; 2438(226)*
g1271 not 2441(240) ; 2441(240)*
g1272 not 2435(225) ; 2435(225)*
g1273 not 2442(239) ; 2442(239)*
g1274 not 2430(224) ; 2430(224)*
g1275 not 2433(242) ; 2433(242)*
g1276 not 2427(223) ; 2427(223)*
g1277 not 2434(241) ; 2434(241)*
g1278 not 2678(232) ; 2678(232)*
g1279 not 2681(351) ; 2681(351)*
g1280 not 2474(231) ; 2474(231)*
g1281 not 2477(369) ; 2477(369)*
g1282 not 2459(325) ; 2459(325)*
g1283 not 2460(326) ; 2460(326)*
g1284 not 1493(327) ; 1493(327)*
g1285 not 1494(328) ; 1494(328)*
g1286 not 1484(329) ; 1484(329)*
g1287 not 1485(330) ; 1485(330)*
g1288 not 1475(331) ; 1475(331)*
g1289 not 1476(332) ; 1476(332)*
g1290 not 2699(248) ; 2699(248)*
g1291 not 2706(340) ; 2706(340)*
g1292 not 2702(250) ; 2702(250)*
g1293 not 2705(339) ; 2705(339)*
g1294 not 2691(252) ; 2691(252)*
g1295 not 2698(344) ; 2698(344)*
g1296 not 2694(254) ; 2694(254)*
g1297 not 2697(342) ; 2697(342)*
g1298 not 2683(256) ; 2683(256)*
g1299 not 2690(348) ; 2690(348)*
g1300 not 2686(258) ; 2686(258)*
g1301 not 2689(346) ; 2689(346)*
g1302 not 2505(266) ; 2505(266)*
g1303 not 2512(355) ; 2512(355)*
g1304 not 2508(268) ; 2508(268)*
g1305 not 2511(353) ; 2511(353)*
g1306 not 2495(270) ; 2495(270)*
g1307 not 2502(359) ; 2502(359)*
g1308 not 2498(272) ; 2498(272)*
g1309 not 2501(357) ; 2501(357)*
g1310 not 2487(274) ; 2487(274)*
g1311 not 2494(363) ; 2494(363)*
g1312 not 2490(276) ; 2490(276)*
g1313 not 2493(361) ; 2493(361)*
g1314 not 2479(278) ; 2479(278)*
g1315 not 2486(367) ; 2486(367)*
g1316 not 2482(280) ; 2482(280)*
g1317 not 2485(365) ; 2485(365)*
g1318 not 2461(285) ; 2461(285)*
g1319 not 2468(373) ; 2468(373)*
g1320 not 2464(287) ; 2464(287)*
g1321 not 2467(371) ; 2467(371)*
g1322 not 1775(416) ; 1775(416)*
g1323 not 1776(323) ; 1776(323)*
g1324 not 1498(417) ; 1498(417)*
g1325 not 1499(324) ; 1499(324)*
g1326 not 2707(428) ; 2707(428)*
g1327 not 2708(427) ; 2708(427)*
g1328 not 1793(432) ; 1793(432)*
g1329 not 1794(430) ; 1794(430)*
g1330 not 1784(436) ; 1784(436)*
g1331 not 1785(434) ; 1785(434)*
g1332 not 2513(441) ; 2513(441)*
g1333 not 2514(439) ; 2514(439)*
g1334 not 2503(445) ; 2503(445)*
g1335 not 2504(443) ; 2504(443)*
g1336 not 1516(449) ; 1516(449)*
g1337 not 1517(447) ; 1517(447)*
g1338 not 1507(453) ; 1507(453)*
g1339 not 1508(451) ; 1508(451)*
g1340 not 2469(458) ; 2469(458)*
g1341 not 2470(456) ; 2470(456)*
g1342 not 2515(553) ; 2515(553)*
g1343 not 2522(539) ; 2522(539)*
g1344 not 2103(247) ; 2103(247)*
g1345 not 1473(545) ; 1473(545)*
g1346 not 2099(249) ; 2099(249)*
g1347 not 1470(562) ; 1470(562)*
g1348 not 2518(418) ; 2518(418)*
g1349 not 2521(595) ; 2521(595)*
g1350 not 2525(549) ; 2525(549)*
g1351 not 2532(590) ; 2532(590)*
g1352 not 2528(550) ; 2528(550)*
g1353 not 2531(589) ; 2531(589)*
g1354 not 560(295) ; 560(295)*
g1355 not 852(619) ; 852(619)*
g1356 not 2631(615) ; 2631(615)*
g1357 not 2638(602) ; 2638(602)*
g1358 not 2523(653) ; 2523(653)*
g1359 not 2524(576) ; 2524(576)*
g1360 not 1540(655) ; 1540(655)*
g1361 not 1541(577) ; 1541(577)*
g1362 not 1537(654) ; 1537(654)*
g1363 not 1538(580) ; 1538(580)*
g1364 not 2665(582) ; 2665(582)*
g1365 not 2672(682) ; 2672(682)*
g1366 not 2778(711) ; 2778(711)*
g1367 not 2781(429) ; 2781(429)*
g1368 not 2770(712) ; 2770(712)*
g1369 not 2773(431) ; 2773(431)*
g1370 not 2762(716) ; 2762(716)*
g1371 not 2765(433) ; 2765(433)*
g1372 not 2754(713) ; 2754(713)*
g1373 not 2757(435) ; 2757(435)*
g1374 not 2746(717) ; 2746(717)*
g1375 not 2749(437) ; 2749(437)*
g1376 not 2738(714) ; 2738(714)*
g1377 not 2741(438) ; 2741(438)*
g1378 not 2533(664) ; 2533(664)*
g1379 not 2534(663) ; 2534(663)*
g1380 not 2626(718) ; 2626(718)*
g1381 not 2629(440) ; 2629(440)*
g1382 not 2618(719) ; 2618(719)*
g1383 not 2621(442) ; 2621(442)*
g1384 not 2610(725) ; 2610(725)*
g1385 not 2613(444) ; 2613(444)*
g1386 not 2602(720) ; 2602(720)*
g1387 not 2605(446) ; 2605(446)*
g1388 not 2594(721) ; 2594(721)*
g1389 not 2597(448) ; 2597(448)*
g1390 not 2586(722) ; 2586(722)*
g1391 not 2589(450) ; 2589(450)*
g1392 not 2578(726) ; 2578(726)*
g1393 not 2581(452) ; 2581(452)*
g1394 not 2570(723) ; 2570(723)*
g1395 not 2573(454) ; 2573(454)*
g1396 not 2562(727) ; 2562(727)*
g1397 not 2565(455) ; 2565(455)*
g1398 not 2554(724) ; 2554(724)*
g1399 not 2557(457) ; 2557(457)*
g1400 not 2634(555) ; 2634(555)*
g1401 not 2637(683) ; 2637(683)*
g1402 not 2642(603) ; 2642(603)*
g1403 not 2645(676) ; 2645(676)*
g1404 not 2639(605) ; 2639(605)*
g1405 not 2646(675) ; 2646(675)*
g1406 not 2650(606) ; 2650(606)*
g1407 not 2653(678) ; 2653(678)*
g1408 not 2647(608) ; 2647(608)*
g1409 not 2654(677) ; 2654(677)*
g1410 not 2658(611) ; 2658(611)*
g1411 not 2661(680) ; 2661(680)*
g1412 not 2655(613) ; 2655(613)*
g1413 not 2662(679) ; 2662(679)*
g1414 not 2668(614) ; 2668(614)*
g1415 not 2671(658) ; 2671(658)*
g1416 not 2151(691) ; 2151(691)*
g1417 not 2158(708) ; 2158(708)*
g1418 not 1820(739) ; 1820(739)*
g1419 not 1821(649) ; 1821(649)*
g1420 not 1823(728) ; 1823(728)*
g1421 not 1824(650) ; 1824(650)*
g1422 not 1543(750) ; 1543(750)*
g1423 not 1544(651) ; 1544(651)*
g1424 not 1546(729) ; 1546(729)*
g1425 not 1547(652) ; 1547(652)*
g1426 not 1542(731) ; 1542(731)*
g1427 not 1539(732) ; 1539(732)*
g1428 not 2673(769) ; 2673(769)*
g1429 not 2674(734) ; 2674(734)*
g1430 not 2775(341) ; 2775(341)*
g1431 not 2782(804) ; 2782(804)*
g1432 not 2767(343) ; 2767(343)*
g1433 not 2774(805) ; 2774(805)*
g1434 not 2759(345) ; 2759(345)*
g1435 not 2766(808) ; 2766(808)*
g1436 not 2751(347) ; 2751(347)*
g1437 not 2758(806) ; 2758(806)*
g1438 not 2743(350) ; 2743(350)*
g1439 not 2750(809) ; 2750(809)*
g1440 not 2735(352) ; 2735(352)*
g1441 not 2742(807) ; 2742(807)*
g1442 not 2623(354) ; 2623(354)*
g1443 not 2630(810) ; 2630(810)*
g1444 not 2615(356) ; 2615(356)*
g1445 not 2622(811) ; 2622(811)*
g1446 not 2607(358) ; 2607(358)*
g1447 not 2614(817) ; 2614(817)*
g1448 not 2599(360) ; 2599(360)*
g1449 not 2606(812) ; 2606(812)*
g1450 not 2591(362) ; 2591(362)*
g1451 not 2598(813) ; 2598(813)*
g1452 not 2583(364) ; 2583(364)*
g1453 not 2590(814) ; 2590(814)*
g1454 not 2575(366) ; 2575(366)*
g1455 not 2582(818) ; 2582(818)*
g1456 not 2567(368) ; 2567(368)*
g1457 not 2574(815) ; 2574(815)*
g1458 not 2559(370) ; 2559(370)*
g1459 not 2566(819) ; 2566(819)*
g1460 not 2551(372) ; 2551(372)*
g1461 not 2558(816) ; 2558(816)*
g1462 not 1752(762) ; 1752(762)*
g1463 not 1753(674) ; 1753(674)*
g1464 not 1761(763) ; 1761(763)*
g1465 not 1762(764) ; 1762(764)*
g1466 not 1770(765) ; 1770(765)*
g1467 not 1771(766) ; 1771(766)*
g1468 not 2663(767) ; 2663(767)*
g1469 not 2664(768) ; 2664(768)*
g1470 not 2110(685) ; 2110(685)*
g1471 not 2113(795) ; 2113(795)*
g1472 not 2164(686) ; 2164(686)*
g1473 not 2167(796) ; 2167(796)*
g1474 not 2115(780) ; 2115(780)*
g1475 not 2122(774) ; 2122(774)*
g1476 not 2169(782) ; 2169(782)*
g1477 not 2176(776) ; 2176(776)*
g1478 not 2126(785) ; 2126(785)*
g1479 not 2129(786) ; 2129(786)*
g1480 not 2107(706) ; 2107(706)*
g1481 not 2114(771) ; 2114(771)*
g1482 not 2161(707) ; 2161(707)*
g1483 not 2168(772) ; 2168(772)*
g1484 not 2154(631) ; 2154(631)*
g1485 not 2157(777) ; 2157(777)*
g1486 not 1825(821) ; 1825(821)*
g1487 not 1822(820) ; 1822(820)*
g1488 not 1548(823) ; 1548(823)*
g1489 not 1545(822) ; 1545(822)*
g1490 not 2535(825) ; 2535(825)*
g1491 not 2542(824) ; 2542(824)*
g1492 not 2059(736) ; 2059(736)*
g1493 not 2060(829) ; 2060(829)*
g1494 not 2055(737) ; 2055(737)*
g1495 not 2056(830) ; 2056(830)*
g1496 not 2051(738) ; 2051(738)*
g1497 not 2052(831) ; 2052(831)*
g1498 not 2047(740) ; 2047(740)*
g1499 not 2048(832) ; 2048(832)*
g1500 not 2043(741) ; 2043(741)*
g1501 not 2044(833) ; 2044(833)*
g1502 not 2039(742) ; 2039(742)*
g1503 not 2040(834) ; 2040(834)*
g1504 not 1597(744) ; 1597(744)*
g1505 not 1598(836) ; 1598(836)*
g1506 not 1593(745) ; 1593(745)*
g1507 not 1594(837) ; 1594(837)*
g1508 not 1589(746) ; 1589(746)*
g1509 not 1590(838) ; 1590(838)*
g1510 not 1585(747) ; 1585(747)*
g1511 not 1586(839) ; 1586(839)*
g1512 not 1581(748) ; 1581(748)*
g1513 not 1582(840) ; 1582(840)*
g1514 not 1577(749) ; 1577(749)*
g1515 not 1578(841) ; 1578(841)*
g1516 not 1573(751) ; 1573(751)*
g1517 not 1574(842) ; 1574(842)*
g1518 not 1569(752) ; 1569(752)*
g1519 not 1570(843) ; 1570(843)*
g1520 not 1565(753) ; 1565(753)*
g1521 not 1566(844) ; 1566(844)*
g1522 not 1561(754) ; 1561(754)*
g1523 not 1562(845) ; 1562(845)*
g1524 not 569(864) ; 569(864)*
g1525 not 570(890) ; 570(890)*
g1526 not 599(865) ; 599(865)*
g1527 not 600(891) ; 600(891)*
g1528 not 2118(688) ; 2118(688)*
g1529 not 2121(869) ; 2121(869)*
g1530 not 2172(690) ; 2172(690)*
g1531 not 2175(871) ; 2175(871)*
g1532 not 2159(892) ; 2159(892)*
g1533 not 2160(778) ; 2160(778)*
g1534 not 2123(697) ; 2123(697)*
g1535 not 2130(875) ; 2130(875)*
g1536 not 2134(787) ; 2134(787)*
g1537 not 2137(882) ; 2137(882)*
g1538 not 2180(788) ; 2180(788)*
g1539 not 2183(883) ; 2183(883)*
g1540 not 2131(789) ; 2131(789)*
g1541 not 2138(880) ; 2138(880)*
g1542 not 2177(790) ; 2177(790)*
g1543 not 2184(881) ; 2184(881)*
g1544 not 2144(791) ; 2144(791)*
g1545 not 2147(888) ; 2147(888)*
g1546 not 2190(792) ; 2190(792)*
g1547 not 2193(889) ; 2193(889)*
g1548 not 2141(793) ; 2141(793)*
g1549 not 2148(884) ; 2148(884)*
g1550 not 2187(794) ; 2187(794)*
g1551 not 2194(885) ; 2194(885)*
g1552 not 2538(730) ; 2538(730)*
g1553 not 2541(902) ; 2541(902)*
g1554 not 2709(827) ; 2709(827)*
g1555 not 2716(928) ; 2716(928)*
g1556 not 2727(899) ; 2727(899)*
g1557 not 2734(584) ; 2734(584)*
g1558 not 2543(900) ; 2543(900)*
g1559 not 2550(835) ; 2550(835)*
g1560 not 2210(933) ; 2210(933)*
g1561 not 2213(852) ; 2213(852)*
g1562 not 2712(861) ; 2712(861)*
g1563 not 2715(904) ; 2715(904)*
g1564 not 578(931) ; 578(931)*
g1565 not 579(866) ; 579(866)*
g1566 not 608(932) ; 608(932)*
g1567 not 609(867) ; 609(867)*
g1568 not 587(874) ; 587(874)*
g1569 not 588(936) ; 588(936)*
g1570 not 2139(939) ; 2139(939)*
g1571 not 2140(943) ; 2140(943)*
g1572 not 2185(940) ; 2185(940)*
g1573 not 2186(944) ; 2186(944)*
g1574 not 2149(947) ; 2149(947)*
g1575 not 2150(949) ; 2150(949)*
g1576 not 2195(948) ; 2195(948)*
g1577 not 2196(950) ; 2196(950)*
g1578 not 1549(963) ; 1549(963)*
g1579 not 1550(901) ; 1550(901)*
g1580 not 2717(1018) ; 2717(1018)*
g1581 not 2718(965) ; 2718(965)*
g1582 not 2730(546) ; 2730(546)*
g1583 not 2733(961) ; 2733(961)*
g1584 not 2546(743) ; 2546(743)*
g1585 not 2549(962) ; 2549(962)*
g1586 not 2207(759) ; 2207(759)*
g1587 not 2214(1025) ; 2214(1025)*
g1588 not 1828(1048) ; 1828(1048)*
g1589 not 1829(966) ; 1829(966)*
g1590 not 1551(1062) ; 1551(1062)*
g1591 not 1552(978) ; 1552(978)*
g1592 not 2215(1009) ; 2215(1009)*
g1593 not 2216(1065) ; 2216(1065)*
g1594 not 1814(1069) ; 1814(1069)*
g1595 not 1815(1010) ; 1815(1010)*
g1596 not 1817(1066) ; 1817(1066)*
g1597 not 1818(1011) ; 1818(1011)*
g1598 not 2200(1031) ; 2200(1031)*
g1599 not 2203(1081) ; 2203(1081)*
g1600 not 2220(1032) ; 2220(1032)*
g1601 not 2223(1082) ; 2223(1082)*
g1602 not 2197(1033) ; 2197(1033)*
g1603 not 2204(1079) ; 2204(1079)*
g1604 not 2217(1034) ; 2217(1034)*
g1605 not 2224(1080) ; 2224(1080)*
g1606 not 1819(1128) ; 1819(1128)*
g1607 not 1816(1127) ; 1816(1127)*
g1608 not 2238(1124) ; 2238(1124)*
g1609 not 2241(770) ; 2241(770)*
g1610 not 2205(1147) ; 2205(1147)*
g1611 not 2206(1149) ; 2206(1149)*
g1612 not 2225(1148) ; 2225(1148)*
g1613 not 2226(1150) ; 2226(1150)*
g1614 not 2719(1190) ; 2719(1190)*
g1615 not 2726(1107) ; 2726(1107)*
g1616 not 635(1189) ; 635(1189)*
g1617 not 636(1125) ; 636(1125)*
g1618 not 638(1188) ; 638(1188)*
g1619 not 639(1126) ; 639(1126)*
g1620 not 2278(1130) ; 2278(1130)*
g1621 not 2281(1212) ; 2281(1212)*
g1622 not 2366(1132) ; 2366(1132)*
g1623 not 2369(1216) ; 2369(1216)*
g1624 not 2270(1134) ; 2270(1134)*
g1625 not 2273(1215) ; 2273(1215)*
g1626 not 2358(1136) ; 2358(1136)*
g1627 not 2361(1219) ; 2361(1219)*
g1628 not 2286(1138) ; 2286(1138)*
g1629 not 2289(1213) ; 2289(1213)*
g1630 not 2374(1140) ; 2374(1140)*
g1631 not 2377(1217) ; 2377(1217)*
g1632 not 2235(684) ; 2235(684)*
g1633 not 2242(1187) ; 2242(1187)*
g1634 not 629(1199) ; 629(1199)*
g1635 not 630(1141) ; 630(1141)*
g1636 not 632(1198) ; 632(1198)*
g1637 not 633(1142) ; 633(1142)*
g1638 not 2347(1185) ; 2347(1185)*
g1639 not 2354(773) ; 2354(773)*
g1640 not 2259(1186) ; 2259(1186)*
g1641 not 2266(775) ; 2266(775)*
g1642 not 2339(1184) ; 2339(1184)*
g1643 not 2346(868) ; 2346(868)*
g1644 not 2251(1183) ; 2251(1183)*
g1645 not 2258(870) ; 2258(870)*
g1646 not 2419(1182) ; 2419(1182)*
g1647 not 2426(872) ; 2426(872)*
g1648 not 2331(1181) ; 2331(1181)*
g1649 not 2338(873) ; 2338(873)*
g1650 not 2294(1152) ; 2294(1152)*
g1651 not 2297(1214) ; 2297(1214)*
g1652 not 2382(1154) ; 2382(1154)*
g1653 not 2385(1218) ; 2385(1218)*
g1654 not 2275(1155) ; 2275(1155)*
g1655 not 2282(1191) ; 2282(1191)*
g1656 not 2283(1156) ; 2283(1156)*
g1657 not 2290(1195) ; 2290(1195)*
g1658 not 2291(1157) ; 2291(1157)*
g1659 not 2298(1208) ; 2298(1208)*
g1660 not 2267(1158) ; 2267(1158)*
g1661 not 2274(1193) ; 2274(1193)*
g1662 not 2363(1159) ; 2363(1159)*
g1663 not 2370(1192) ; 2370(1192)*
g1664 not 2371(1160) ; 2371(1160)*
g1665 not 2378(1196) ; 2378(1196)*
g1666 not 2379(1161) ; 2379(1161)*
g1667 not 2386(1209) ; 2386(1209)*
g1668 not 2355(1162) ; 2355(1162)*
g1669 not 2362(1194) ; 2362(1194)*
g1670 not 2299(1164) ; 2299(1164)*
g1671 not 2306(1233) ; 2306(1233)*
g1672 not 2307(1166) ; 2307(1166)*
g1673 not 2314(1232) ; 2314(1232)*
g1674 not 2387(1168) ; 2387(1168)*
g1675 not 2394(1237) ; 2394(1237)*
g1676 not 2395(1170) ; 2395(1170)*
g1677 not 2402(1236) ; 2402(1236)*
g1678 not 2310(1173) ; 2310(1173)*
g1679 not 2313(1223) ; 2313(1223)*
g1680 not 2302(1174) ; 2302(1174)*
g1681 not 2305(1222) ; 2305(1222)*
g1682 not 2398(1177) ; 2398(1177)*
g1683 not 2401(1227) ; 2401(1227)*
g1684 not 2390(1178) ; 2390(1178)*
g1685 not 2393(1226) ; 2393(1226)*
g1686 not 2722(1047) ; 2722(1047)*
g1687 not 2725(1247) ; 2725(1247)*
g1688 not 640(1246) ; 640(1246)*
g1689 not 637(1245) ; 637(1245)*
g1690 not 908(1248) ; 908(1248)*
g1691 not 909(1267) ; 909(1267)*
g1692 not 1126(1249) ; 1126(1249)*
g1693 not 1127(1271) ; 1127(1271)*
g1694 not 899(1250) ; 899(1250)*
g1695 not 900(1270) ; 900(1270)*
g1696 not 1117(1251) ; 1117(1251)*
g1697 not 1118(1274) ; 1118(1274)*
g1698 not 916(1252) ; 916(1252)*
g1699 not 917(1268) ; 917(1268)*
g1700 not 1134(1253) ; 1134(1253)*
g1701 not 1135(1272) ; 1135(1272)*
g1702 not 645(1197) ; 645(1197)*
g1703 not 646(1254) ; 646(1254)*
g1704 not 634(1256) ; 634(1256)*
g1705 not 631(1255) ; 631(1255)*
g1706 not 2350(687) ; 2350(687)*
g1707 not 2353(1243) ; 2353(1243)*
g1708 not 2262(689) ; 2262(689)*
g1709 not 2265(1244) ; 2265(1244)*
g1710 not 2342(779) ; 2342(779)*
g1711 not 2345(1242) ; 2345(1242)*
g1712 not 2254(781) ; 2254(781)*
g1713 not 2257(1241) ; 2257(1241)*
g1714 not 2422(783) ; 2422(783)*
g1715 not 2425(1240) ; 2425(1240)*
g1716 not 2334(784) ; 2334(784)*
g1717 not 2337(1239) ; 2337(1239)*
g1718 not 925(1265) ; 925(1265)*
g1719 not 926(1269) ; 926(1269)*
g1720 not 1143(1266) ; 1143(1266)*
g1721 not 1144(1273) ; 1144(1273)*
g1722 not 928(1292) ; 928(1292)*
g1723 not 929(1279) ; 929(1279)*
g1724 not 938(1291) ; 938(1291)*
g1725 not 939(1280) ; 939(1280)*
g1726 not 2315(1281) ; 2315(1281)*
g1727 not 2322(1290) ; 2322(1290)*
g1728 not 2323(1282) ; 2323(1282)*
g1729 not 2330(1287) ; 2330(1287)*
g1730 not 1146(1298) ; 1146(1298)*
g1731 not 1147(1283) ; 1147(1283)*
g1732 not 1156(1297) ; 1156(1297)*
g1733 not 1157(1284) ; 1157(1284)*
g1734 not 2403(1285) ; 2403(1285)*
g1735 not 2410(1296) ; 2410(1296)*
g1736 not 2411(1286) ; 2411(1286)*
g1737 not 2418(1293) ; 2418(1293)*
g1738 not 1826(1299) ; 1826(1299)*
g1739 not 1827(1238) ; 1827(1238)*
g1740 not 1114(1309) ; 1114(1309)*
g1741 not 1115(1257) ; 1115(1257)*
g1742 not 683(1310) ; 683(1310)*
g1743 not 684(1258) ; 684(1258)*
g1744 not 1098(1311) ; 1098(1311)*
g1745 not 1099(1259) ; 1099(1259)*
g1746 not 664(1312) ; 664(1312)*
g1747 not 665(1260) ; 665(1260)*
g1748 not 1180(1313) ; 1180(1313)*
g1749 not 1181(1261) ; 1181(1261)*
g1750 not 962(1314) ; 962(1314)*
g1751 not 963(1262) ; 963(1262)*
g1752 not 2227(1308) ; 2227(1308)*
g1753 not 2234(1263) ; 2234(1263)*
g1754 not 2243(1300) ; 2243(1300)*
g1755 not 2250(1264) ; 2250(1264)*
g1756 not 2326(1230) ; 2326(1230)*
g1757 not 2329(1322) ; 2329(1322)*
g1758 not 2318(1231) ; 2318(1231)*
g1759 not 2321(1320) ; 2321(1320)*
g1760 not 2414(1234) ; 2414(1234)*
g1761 not 2417(1328) ; 2417(1328)*
g1762 not 2406(1235) ; 2406(1235)*
g1763 not 2409(1326) ; 2409(1326)*
g1764 not 2230(1206) ; 2230(1206)*
g1765 not 2233(1338) ; 2233(1338)*
g1766 not 2246(1207) ; 2246(1207)*
g1767 not 2249(1331) ; 2249(1331)*
g1768 not 947(1353) ; 947(1353)*
g1769 not 948(1319) ; 948(1319)*
g1770 not 955(1351) ; 955(1351)*
g1771 not 956(1321) ; 956(1321)*
g1772 not 1165(1356) ; 1165(1356)*
g1773 not 1166(1325) ; 1166(1325)*
g1774 not 1173(1354) ; 1173(1354)*
g1775 not 1174(1327) ; 1174(1327)*
g1776 not 641(1365) ; 641(1365)*
g1777 not 642(1345) ; 642(1345)*
g1778 not 648(1366) ; 648(1366)*
g1779 not 649(1346) ; 649(1346)*
g1780 not 976(1373) ; 976(1373)*
g1781 not 969(1359) ; 969(1359)*
g1782 not 1193(1374) ; 1193(1374)*
g1783 not 1186(1360) ; 1186(1360)*
g1784 not 329(1414) ; 329(1414)*
g1785 not 991(1411) ; 991(1411)*
