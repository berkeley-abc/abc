name C1355.iscas
i 1GAT(0)
i 8GAT(1)
i 15GAT(2)
i 22GAT(3)
i 29GAT(4)
i 36GAT(5)
i 43GAT(6)
i 50GAT(7)
i 57GAT(8)
i 64GAT(9)
i 71GAT(10)
i 78GAT(11)
i 85GAT(12)
i 92GAT(13)
i 99GAT(14)
i 106GAT(15)
i 113GAT(16)
i 120GAT(17)
i 127GAT(18)
i 134GAT(19)
i 141GAT(20)
i 148GAT(21)
i 155GAT(22)
i 162GAT(23)
i 169GAT(24)
i 176GAT(25)
i 183GAT(26)
i 190GAT(27)
i 197GAT(28)
i 204GAT(29)
i 211GAT(30)
i 218GAT(31)
i 225GAT(32)
i 226GAT(33)
i 227GAT(34)
i 228GAT(35)
i 229GAT(36)
i 230GAT(37)
i 231GAT(38)
i 232GAT(39)
i 233GAT(40)

o 1324GAT(583)
o 1325GAT(579)
o 1326GAT(575)
o 1327GAT(571)
o 1328GAT(584)
o 1329GAT(580)
o 1330GAT(576)
o 1331GAT(572)
o 1332GAT(585)
o 1333GAT(581)
o 1334GAT(577)
o 1335GAT(573)
o 1336GAT(586)
o 1337GAT(582)
o 1338GAT(578)
o 1339GAT(574)
o 1340GAT(567)
o 1341GAT(563)
o 1342GAT(559)
o 1343GAT(555)
o 1344GAT(568)
o 1345GAT(564)
o 1346GAT(560)
o 1347GAT(556)
o 1348GAT(569)
o 1349GAT(565)
o 1350GAT(561)
o 1351GAT(557)
o 1352GAT(570)
o 1353GAT(566)
o 1354GAT(562)
o 1355GAT(558)

g1 and 233GAT(40) 232GAT(39) ; 263GAT(41)
g2 and 233GAT(40) 231GAT(38) ; 260GAT(42)
g3 and 233GAT(40) 230GAT(37) ; 257GAT(43)
g4 and 233GAT(40) 229GAT(36) ; 254GAT(44)
g5 and 233GAT(40) 228GAT(35) ; 251GAT(45)
g6 and 233GAT(40) 227GAT(34) ; 248GAT(46)
g7 and 233GAT(40) 226GAT(33) ; 245GAT(47)
g8 and 233GAT(40) 225GAT(32) ; 242GAT(48)
g9 and 218GAT(31) 211GAT(30) ; 311GAT(49)
g10 and 204GAT(29) 197GAT(28) ; 308GAT(50)
g11 and 218GAT(31) 190GAT(27) ; 359GAT(51)
g12 and 211GAT(30) 183GAT(26) ; 353GAT(52)
g13 and 190GAT(27) 183GAT(26) ; 305GAT(53)
g14 and 204GAT(29) 176GAT(25) ; 347GAT(54)
g15 and 197GAT(28) 169GAT(24) ; 341GAT(55)
g16 and 176GAT(25) 169GAT(24) ; 302GAT(56)
g17 and 162GAT(23) 155GAT(22) ; 299GAT(57)
g18 and 148GAT(21) 141GAT(20) ; 296GAT(58)
g19 and 162GAT(23) 134GAT(19) ; 356GAT(59)
g20 and 155GAT(22) 127GAT(18) ; 350GAT(60)
g21 and 134GAT(19) 127GAT(18) ; 293GAT(61)
g22 and 148GAT(21) 120GAT(17) ; 344GAT(62)
g23 and 141GAT(20) 113GAT(16) ; 338GAT(63)
g24 and 120GAT(17) 113GAT(16) ; 290GAT(64)
g25 and 106GAT(15) 99GAT(14) ; 287GAT(65)
g26 and 92GAT(13) 85GAT(12) ; 284GAT(66)
g27 and 106GAT(15) 78GAT(11) ; 335GAT(67)
g28 and 99GAT(14) 71GAT(10) ; 329GAT(68)
g29 and 78GAT(11) 71GAT(10) ; 281GAT(69)
g30 and 92GAT(13) 64GAT(9) ; 323GAT(70)
g31 and 85GAT(12) 57GAT(8) ; 317GAT(71)
g32 and 64GAT(9) 57GAT(8) ; 278GAT(72)
g33 and 50GAT(7) 43GAT(6) ; 275GAT(73)
g34 and 36GAT(5) 29GAT(4) ; 272GAT(74)
g35 and 50GAT(7) 22GAT(3) ; 332GAT(75)
g36 and 43GAT(6) 15GAT(2) ; 326GAT(76)
g37 and 22GAT(3) 15GAT(2) ; 269GAT(77)
g38 and 36GAT(5) 8GAT(1) ; 320GAT(78)
g39 and 29GAT(4) 1GAT(0) ; 314GAT(79)
g40 and 8GAT(1) 1GAT(0) ; 266GAT(80)
g41 and 359GAT(51) 218GAT(31) ; 425GAT(81)
g42 and 311GAT(49) 218GAT(31) ; 393GAT(82)
g43 and 353GAT(52) 211GAT(30) ; 421GAT(83)
g44 and 311GAT(49) 211GAT(30) ; 392GAT(84)
g45 and 347GAT(54) 204GAT(29) ; 417GAT(85)
g46 and 308GAT(50) 204GAT(29) ; 391GAT(86)
g47 and 341GAT(55) 197GAT(28) ; 413GAT(87)
g48 and 308GAT(50) 197GAT(28) ; 390GAT(88)
g49 and 359GAT(51) 190GAT(27) ; 424GAT(89)
g50 and 305GAT(53) 190GAT(27) ; 389GAT(90)
g51 and 353GAT(52) 183GAT(26) ; 420GAT(91)
g52 and 305GAT(53) 183GAT(26) ; 388GAT(92)
g53 and 347GAT(54) 176GAT(25) ; 416GAT(93)
g54 and 302GAT(56) 176GAT(25) ; 387GAT(94)
g55 and 341GAT(55) 169GAT(24) ; 412GAT(95)
g56 and 302GAT(56) 169GAT(24) ; 386GAT(96)
g57 and 356GAT(59) 162GAT(23) ; 423GAT(97)
g58 and 299GAT(57) 162GAT(23) ; 385GAT(98)
g59 and 350GAT(60) 155GAT(22) ; 419GAT(99)
g60 and 299GAT(57) 155GAT(22) ; 384GAT(100)
g61 and 344GAT(62) 148GAT(21) ; 415GAT(101)
g62 and 296GAT(58) 148GAT(21) ; 383GAT(102)
g63 and 338GAT(63) 141GAT(20) ; 411GAT(103)
g64 and 296GAT(58) 141GAT(20) ; 382GAT(104)
g65 and 356GAT(59) 134GAT(19) ; 422GAT(105)
g66 and 293GAT(61) 134GAT(19) ; 381GAT(106)
g67 and 350GAT(60) 127GAT(18) ; 418GAT(107)
g68 and 293GAT(61) 127GAT(18) ; 380GAT(108)
g69 and 344GAT(62) 120GAT(17) ; 414GAT(109)
g70 and 290GAT(64) 120GAT(17) ; 379GAT(110)
g71 and 338GAT(63) 113GAT(16) ; 410GAT(111)
g72 and 290GAT(64) 113GAT(16) ; 378GAT(112)
g73 and 335GAT(67) 106GAT(15) ; 409GAT(113)
g74 and 287GAT(65) 106GAT(15) ; 377GAT(114)
g75 and 329GAT(68) 99GAT(14) ; 405GAT(115)
g76 and 287GAT(65) 99GAT(14) ; 376GAT(116)
g77 and 323GAT(70) 92GAT(13) ; 401GAT(117)
g78 and 284GAT(66) 92GAT(13) ; 375GAT(118)
g79 and 317GAT(71) 85GAT(12) ; 397GAT(119)
g80 and 284GAT(66) 85GAT(12) ; 374GAT(120)
g81 and 335GAT(67) 78GAT(11) ; 408GAT(121)
g82 and 281GAT(69) 78GAT(11) ; 373GAT(122)
g83 and 329GAT(68) 71GAT(10) ; 404GAT(123)
g84 and 281GAT(69) 71GAT(10) ; 372GAT(124)
g85 and 323GAT(70) 64GAT(9) ; 400GAT(125)
g86 and 278GAT(72) 64GAT(9) ; 371GAT(126)
g87 and 317GAT(71) 57GAT(8) ; 396GAT(127)
g88 and 278GAT(72) 57GAT(8) ; 370GAT(128)
g89 and 332GAT(75) 50GAT(7) ; 407GAT(129)
g90 and 275GAT(73) 50GAT(7) ; 369GAT(130)
g91 and 326GAT(76) 43GAT(6) ; 403GAT(131)
g92 and 275GAT(73) 43GAT(6) ; 368GAT(132)
g93 and 320GAT(78) 36GAT(5) ; 399GAT(133)
g94 and 272GAT(74) 36GAT(5) ; 367GAT(134)
g95 and 314GAT(79) 29GAT(4) ; 395GAT(135)
g96 and 272GAT(74) 29GAT(4) ; 366GAT(136)
g97 and 332GAT(75) 22GAT(3) ; 406GAT(137)
g98 and 269GAT(77) 22GAT(3) ; 365GAT(138)
g99 and 326GAT(76) 15GAT(2) ; 402GAT(139)
g100 and 269GAT(77) 15GAT(2) ; 364GAT(140)
g101 and 320GAT(78) 8GAT(1) ; 398GAT(141)
g102 and 266GAT(80) 8GAT(1) ; 363GAT(142)
g103 and 314GAT(79) 1GAT(0) ; 394GAT(143)
g104 and 266GAT(80) 1GAT(0) ; 362GAT(144)
g105 and 425GAT(81) 424GAT(89) ; 519GAT(145)
g106 and 393GAT(82) 392GAT(84) ; 471GAT(146)
g107 and 421GAT(83) 420GAT(91) ; 513GAT(147)
g108 and 417GAT(85) 416GAT(93) ; 507GAT(148)
g109 and 391GAT(86) 390GAT(88) ; 468GAT(149)
g110 and 413GAT(87) 412GAT(95) ; 501GAT(150)
g111 and 389GAT(90) 388GAT(92) ; 465GAT(151)
g112 and 387GAT(94) 386GAT(96) ; 462GAT(152)
g113 and 423GAT(97) 422GAT(105) ; 516GAT(153)
g114 and 385GAT(98) 384GAT(100) ; 459GAT(154)
g115 and 419GAT(99) 418GAT(107) ; 510GAT(155)
g116 and 415GAT(101) 414GAT(109) ; 504GAT(156)
g117 and 383GAT(102) 382GAT(104) ; 456GAT(157)
g118 and 411GAT(103) 410GAT(111) ; 498GAT(158)
g119 and 381GAT(106) 380GAT(108) ; 453GAT(159)
g120 and 379GAT(110) 378GAT(112) ; 450GAT(160)
g121 and 409GAT(113) 408GAT(121) ; 495GAT(161)
g122 and 377GAT(114) 376GAT(116) ; 447GAT(162)
g123 and 405GAT(115) 404GAT(123) ; 489GAT(163)
g124 and 401GAT(117) 400GAT(125) ; 483GAT(164)
g125 and 375GAT(118) 374GAT(120) ; 444GAT(165)
g126 and 397GAT(119) 396GAT(127) ; 477GAT(166)
g127 and 373GAT(122) 372GAT(124) ; 441GAT(167)
g128 and 371GAT(126) 370GAT(128) ; 438GAT(168)
g129 and 407GAT(129) 406GAT(137) ; 492GAT(169)
g130 and 369GAT(130) 368GAT(132) ; 435GAT(170)
g131 and 403GAT(131) 402GAT(139) ; 486GAT(171)
g132 and 399GAT(133) 398GAT(141) ; 480GAT(172)
g133 and 367GAT(134) 366GAT(136) ; 432GAT(173)
g134 and 395GAT(135) 394GAT(143) ; 474GAT(174)
g135 and 365GAT(138) 364GAT(140) ; 429GAT(175)
g136 and 363GAT(142) 362GAT(144) ; 426GAT(176)
g137 and 519GAT(145) 516GAT(153) ; 567GAT(177)
g138 and 471GAT(146) 468GAT(149) ; 543GAT(178)
g139 and 513GAT(147) 510GAT(155) ; 564GAT(179)
g140 and 507GAT(148) 504GAT(156) ; 561GAT(180)
g141 and 501GAT(150) 498GAT(158) ; 558GAT(181)
g142 and 465GAT(151) 462GAT(152) ; 540GAT(182)
g143 and 459GAT(154) 456GAT(157) ; 537GAT(183)
g144 and 453GAT(159) 450GAT(160) ; 534GAT(184)
g145 and 495GAT(161) 492GAT(169) ; 555GAT(185)
g146 and 447GAT(162) 444GAT(165) ; 531GAT(186)
g147 and 489GAT(163) 486GAT(171) ; 552GAT(187)
g148 and 483GAT(164) 480GAT(172) ; 549GAT(188)
g149 and 477GAT(166) 474GAT(174) ; 546GAT(189)
g150 and 441GAT(167) 438GAT(168) ; 528GAT(190)
g151 and 435GAT(170) 432GAT(173) ; 525GAT(191)
g152 and 429GAT(175) 426GAT(176) ; 522GAT(192)
g153 and 567GAT(177) 519GAT(145) ; 601GAT(193)
g154 and 543GAT(178) 471GAT(146) ; 585GAT(194)
g155 and 564GAT(179) 513GAT(147) ; 599GAT(195)
g156 and 561GAT(180) 507GAT(148) ; 597GAT(196)
g157 and 543GAT(178) 468GAT(149) ; 584GAT(197)
g158 and 558GAT(181) 501GAT(150) ; 595GAT(198)
g159 and 540GAT(182) 465GAT(151) ; 583GAT(199)
g160 and 540GAT(182) 462GAT(152) ; 582GAT(200)
g161 and 567GAT(177) 516GAT(153) ; 600GAT(201)
g162 and 537GAT(183) 459GAT(154) ; 581GAT(202)
g163 and 564GAT(179) 510GAT(155) ; 598GAT(203)
g164 and 561GAT(180) 504GAT(156) ; 596GAT(204)
g165 and 537GAT(183) 456GAT(157) ; 580GAT(205)
g166 and 558GAT(181) 498GAT(158) ; 594GAT(206)
g167 and 534GAT(184) 453GAT(159) ; 579GAT(207)
g168 and 534GAT(184) 450GAT(160) ; 578GAT(208)
g169 and 555GAT(185) 495GAT(161) ; 593GAT(209)
g170 and 531GAT(186) 447GAT(162) ; 577GAT(210)
g171 and 552GAT(187) 489GAT(163) ; 591GAT(211)
g172 and 549GAT(188) 483GAT(164) ; 589GAT(212)
g173 and 531GAT(186) 444GAT(165) ; 576GAT(213)
g174 and 546GAT(189) 477GAT(166) ; 587GAT(214)
g175 and 528GAT(190) 441GAT(167) ; 575GAT(215)
g176 and 528GAT(190) 438GAT(168) ; 574GAT(216)
g177 and 555GAT(185) 492GAT(169) ; 592GAT(217)
g178 and 525GAT(191) 435GAT(170) ; 573GAT(218)
g179 and 552GAT(187) 486GAT(171) ; 590GAT(219)
g180 and 549GAT(188) 480GAT(172) ; 588GAT(220)
g181 and 525GAT(191) 432GAT(173) ; 572GAT(221)
g182 and 546GAT(189) 474GAT(174) ; 586GAT(222)
g183 and 522GAT(192) 429GAT(175) ; 571GAT(223)
g184 and 522GAT(192) 426GAT(176) ; 570GAT(224)
g185 and 601GAT(193) 600GAT(201) ; 663GAT(225)
g186 and 585GAT(194) 584GAT(197) ; 637GAT(226)
g187 and 599GAT(195) 598GAT(203) ; 660GAT(227)
g188 and 597GAT(196) 596GAT(204) ; 657GAT(228)
g189 and 595GAT(198) 594GAT(206) ; 654GAT(229)
g190 and 583GAT(199) 582GAT(200) ; 632GAT(230)
g191 and 581GAT(202) 580GAT(205) ; 627GAT(231)
g192 and 579GAT(207) 578GAT(208) ; 622GAT(232)
g193 and 593GAT(209) 592GAT(217) ; 651GAT(233)
g194 and 577GAT(210) 576GAT(213) ; 617GAT(234)
g195 and 591GAT(211) 590GAT(219) ; 648GAT(235)
g196 and 589GAT(212) 588GAT(220) ; 645GAT(236)
g197 and 587GAT(214) 586GAT(222) ; 642GAT(237)
g198 and 575GAT(215) 574GAT(216) ; 612GAT(238)
g199 and 573GAT(218) 572GAT(221) ; 607GAT(239)
g200 and 571GAT(223) 570GAT(224) ; 602GAT(240)
g201 and 637GAT(226) 632GAT(230) ; 681GAT(241)
g202 and 637GAT(226) 627GAT(231) ; 687GAT(242)
g203 and 632GAT(230) 622GAT(232) ; 684GAT(243)
g204 and 627GAT(231) 622GAT(232) ; 678GAT(244)
g205 and 617GAT(234) 612GAT(238) ; 669GAT(245)
g206 and 617GAT(234) 607GAT(239) ; 675GAT(246)
g207 and 612GAT(238) 602GAT(240) ; 672GAT(247)
g208 and 607GAT(239) 602GAT(240) ; 666GAT(248)
g209 and 681GAT(241) 637GAT(226) ; 701GAT(249)
g210 and 687GAT(242) 637GAT(226) ; 705GAT(250)
g211 and 681GAT(241) 632GAT(230) ; 700GAT(251)
g212 and 684GAT(243) 632GAT(230) ; 703GAT(252)
g213 and 678GAT(244) 627GAT(231) ; 699GAT(253)
g214 and 687GAT(242) 627GAT(231) ; 704GAT(254)
g215 and 678GAT(244) 622GAT(232) ; 698GAT(255)
g216 and 684GAT(243) 622GAT(232) ; 702GAT(256)
g217 and 669GAT(245) 617GAT(234) ; 693GAT(257)
g218 and 675GAT(246) 617GAT(234) ; 697GAT(258)
g219 and 669GAT(245) 612GAT(238) ; 692GAT(259)
g220 and 672GAT(247) 612GAT(238) ; 695GAT(260)
g221 and 666GAT(248) 607GAT(239) ; 691GAT(261)
g222 and 675GAT(246) 607GAT(239) ; 696GAT(262)
g223 and 666GAT(248) 602GAT(240) ; 690GAT(263)
g224 and 672GAT(247) 602GAT(240) ; 694GAT(264)
g225 and 701GAT(249) 700GAT(251) ; 721GAT(265)
g226 and 705GAT(250) 704GAT(254) ; 727GAT(266)
g227 and 703GAT(252) 702GAT(256) ; 724GAT(267)
g228 and 699GAT(253) 698GAT(255) ; 718GAT(268)
g229 and 693GAT(257) 692GAT(259) ; 709GAT(269)
g230 and 697GAT(258) 696GAT(262) ; 715GAT(270)
g231 and 695GAT(260) 694GAT(264) ; 712GAT(271)
g232 and 691GAT(261) 690GAT(263) ; 706GAT(272)
g233 and 715GAT(270) 263GAT(41) ; 751GAT(273)
g234 and 712GAT(271) 260GAT(42) ; 748GAT(274)
g235 and 709GAT(269) 257GAT(43) ; 745GAT(275)
g236 and 706GAT(272) 254GAT(44) ; 742GAT(276)
g237 and 727GAT(266) 251GAT(45) ; 739GAT(277)
g238 and 724GAT(267) 248GAT(46) ; 736GAT(278)
g239 and 721GAT(265) 245GAT(47) ; 733GAT(279)
g240 and 718GAT(268) 242GAT(48) ; 730GAT(280)
g241 and 751GAT(273) 263GAT(41) ; 768GAT(281)
g242 and 748GAT(274) 260GAT(42) ; 766GAT(282)
g243 and 745GAT(275) 257GAT(43) ; 764GAT(283)
g244 and 742GAT(276) 254GAT(44) ; 762GAT(284)
g245 and 739GAT(277) 251GAT(45) ; 760GAT(285)
g246 and 736GAT(278) 248GAT(46) ; 758GAT(286)
g247 and 733GAT(279) 245GAT(47) ; 756GAT(287)
g248 and 730GAT(280) 242GAT(48) ; 754GAT(288)
g249 and 733GAT(279) 721GAT(265) ; 757GAT(289)
g250 and 739GAT(277) 727GAT(266) ; 761GAT(290)
g251 and 736GAT(278) 724GAT(267) ; 759GAT(291)
g252 and 730GAT(280) 718GAT(268) ; 755GAT(292)
g253 and 745GAT(275) 709GAT(269) ; 765GAT(293)
g254 and 751GAT(273) 715GAT(270) ; 769GAT(294)
g255 and 748GAT(274) 712GAT(271) ; 767GAT(295)
g256 and 742GAT(276) 706GAT(272) ; 763GAT(296)
g257 and 769GAT(294) 768GAT(281) ; 791GAT(297)
g258 and 767GAT(295) 766GAT(282) ; 788GAT(298)
g259 and 765GAT(293) 764GAT(283) ; 785GAT(299)
g260 and 763GAT(296) 762GAT(284) ; 782GAT(300)
g261 and 761GAT(290) 760GAT(285) ; 779GAT(301)
g262 and 759GAT(291) 758GAT(286) ; 776GAT(302)
g263 and 757GAT(289) 756GAT(287) ; 773GAT(303)
g264 and 755GAT(292) 754GAT(288) ; 770GAT(304)
g265 and 791GAT(297) 663GAT(225) ; 815GAT(305)
g266 and 788GAT(298) 660GAT(227) ; 812GAT(306)
g267 and 785GAT(299) 657GAT(228) ; 809GAT(307)
g268 and 782GAT(300) 654GAT(229) ; 806GAT(308)
g269 and 779GAT(301) 651GAT(233) ; 803GAT(309)
g270 and 776GAT(302) 648GAT(235) ; 800GAT(310)
g271 and 773GAT(303) 645GAT(236) ; 797GAT(311)
g272 and 770GAT(304) 642GAT(237) ; 794GAT(312)
g273 and 815GAT(305) 791GAT(297) ; 833GAT(313)
g274 and 812GAT(306) 788GAT(298) ; 831GAT(314)
g275 and 809GAT(307) 785GAT(299) ; 829GAT(315)
g276 and 806GAT(308) 782GAT(300) ; 827GAT(316)
g277 and 803GAT(309) 779GAT(301) ; 825GAT(317)
g278 and 800GAT(310) 776GAT(302) ; 823GAT(318)
g279 and 797GAT(311) 773GAT(303) ; 821GAT(319)
g280 and 794GAT(312) 770GAT(304) ; 819GAT(320)
g281 and 815GAT(305) 663GAT(225) ; 832GAT(321)
g282 and 812GAT(306) 660GAT(227) ; 830GAT(322)
g283 and 809GAT(307) 657GAT(228) ; 828GAT(323)
g284 and 806GAT(308) 654GAT(229) ; 826GAT(324)
g285 and 803GAT(309) 651GAT(233) ; 824GAT(325)
g286 and 800GAT(310) 648GAT(235) ; 822GAT(326)
g287 and 797GAT(311) 645GAT(236) ; 820GAT(327)
g288 and 794GAT(312) 642GAT(237) ; 818GAT(328)
g289 and 833GAT(313) 832GAT(321) ; 899GAT(329)
g290 and 831GAT(314) 830GAT(322) ; 912GAT(330)
g291 and 829GAT(315) 828GAT(323) ; 886GAT(331)
g292 and 827GAT(316) 826GAT(324) ; 925GAT(332)
g293 and 825GAT(317) 824GAT(325) ; 873GAT(333)
g294 and 823GAT(318) 822GAT(326) ; 860GAT(334)
g295 and 821GAT(319) 820GAT(327) ; 847GAT(335)
g296 and 819GAT(320) 818GAT(328) ; 834GAT(336)
g297 and 899GAT(329) ; 951GAT(337)
g298 and 899GAT(329) ; 955GAT(338)
g299 and 899GAT(329) ; 963GAT(339)
g300 and 899GAT(329) ; 966GAT(340)
g301 and 899GAT(329) ; 969GAT(341)
g302 and 912GAT(330) ; 953GAT(342)
g303 and 912GAT(330) ; 957GAT(343)
g304 and 912GAT(330) ; 960GAT(344)
g305 and 912GAT(330) ; 965GAT(345)
g306 and 912GAT(330) ; 968GAT(346)
g307 and 886GAT(331) ; 950GAT(347)
g308 and 886GAT(331) ; 952GAT(348)
g309 and 886GAT(331) ; 959GAT(349)
g310 and 886GAT(331) ; 962GAT(350)
g311 and 886GAT(331) ; 967GAT(351)
g312 and 925GAT(332) ; 954GAT(352)
g313 and 925GAT(332) ; 956GAT(353)
g314 and 925GAT(332) ; 958GAT(354)
g315 and 925GAT(332) ; 961GAT(355)
g316 and 925GAT(332) ; 964GAT(356)
g317 and 873GAT(333) ; 943GAT(357)
g318 and 873GAT(333) ; 946GAT(358)
g319 and 873GAT(333) ; 949GAT(359)
g320 and 873GAT(333) ; 971GAT(360)
g321 and 873GAT(333) ; 975GAT(361)
g322 and 860GAT(334) ; 940GAT(362)
g323 and 860GAT(334) ; 945GAT(363)
g324 and 860GAT(334) ; 948GAT(364)
g325 and 860GAT(334) ; 973GAT(365)
g326 and 860GAT(334) ; 977GAT(366)
g327 and 847GAT(335) ; 939GAT(367)
g328 and 847GAT(335) ; 942GAT(368)
g329 and 847GAT(335) ; 947GAT(369)
g330 and 847GAT(335) ; 970GAT(370)
g331 and 847GAT(335) ; 972GAT(371)
g332 and 834GAT(336) ; 938GAT(372)
g333 and 834GAT(336) ; 941GAT(373)
g334 and 834GAT(336) ; 944GAT(374)
g335 and 834GAT(336) ; 974GAT(375)
g336 and 834GAT(336) ; 976GAT(376)
g337 and 899GAT(329) 960GAT(344) 959GAT(349) 958GAT(354) ; 982GAT(377)
g338 and 963GAT(339) 912GAT(330) 962GAT(350) 961GAT(355) ; 983GAT(378)
g339 and 966GAT(340) 965GAT(345) 886GAT(331) 964GAT(356) ; 984GAT(379)
g340 and 969GAT(341) 968GAT(346) 967GAT(351) 925GAT(332) ; 985GAT(380)
g341 and 873GAT(333) 940GAT(362) 939GAT(367) 938GAT(372) ; 978GAT(381)
g342 and 943GAT(357) 860GAT(334) 942GAT(368) 941GAT(373) ; 979GAT(382)
g343 and 946GAT(358) 945GAT(363) 847GAT(335) 944GAT(374) ; 980GAT(383)
g344 and 949GAT(359) 948GAT(364) 947GAT(369) 834GAT(336) ; 981GAT(384)
g345 and 985GAT(380)* 984GAT(379)* 983GAT(378)* 982GAT(377)* ; 991GAT(385)
g346 and 981GAT(384)* 980GAT(383)* 979GAT(382)* 978GAT(381)* ; 986GAT(386)
g347 and 986GAT(386) 899GAT(329) 953GAT(342) 952GAT(348) 925GAT(332) ; 1001GAT(387)
g348 and 986GAT(386) 899GAT(329) 957GAT(343) 886GAT(331) 956GAT(353) ; 1011GAT(388)
g349 and 986GAT(386) 951GAT(337) 912GAT(330) 950GAT(347) 925GAT(332) ; 996GAT(389)
g350 and 986GAT(386) 955GAT(338) 912GAT(330) 886GAT(331) 954GAT(352) ; 1006GAT(390)
g351 and 991GAT(385) 873GAT(333) 973GAT(365) 972GAT(371) 834GAT(336) ; 1021GAT(391)
g352 and 991GAT(385) 873GAT(333) 977GAT(366) 847GAT(335) 976GAT(376) ; 1031GAT(392)
g353 and 991GAT(385) 971GAT(360) 860GAT(334) 970GAT(370) 834GAT(336) ; 1016GAT(393)
g354 and 991GAT(385) 975GAT(361) 860GAT(334) 847GAT(335) 974GAT(375) ; 1026GAT(394)
g355 and 1016GAT(393) 899GAT(329) ; 1093GAT(395)
g356 and 1021GAT(391) 899GAT(329) ; 1105GAT(396)
g357 and 1026GAT(394) 899GAT(329) ; 1117GAT(397)
g358 and 1031GAT(392) 899GAT(329) ; 1129GAT(398)
g359 and 1016GAT(393) 912GAT(330) ; 1090GAT(399)
g360 and 1021GAT(391) 912GAT(330) ; 1102GAT(400)
g361 and 1026GAT(394) 912GAT(330) ; 1114GAT(401)
g362 and 1031GAT(392) 912GAT(330) ; 1126GAT(402)
g363 and 1016GAT(393) 886GAT(331) ; 1087GAT(403)
g364 and 1021GAT(391) 886GAT(331) ; 1099GAT(404)
g365 and 1026GAT(394) 886GAT(331) ; 1111GAT(405)
g366 and 1031GAT(392) 886GAT(331) ; 1123GAT(406)
g367 and 1016GAT(393) 925GAT(332) ; 1084GAT(407)
g368 and 1021GAT(391) 925GAT(332) ; 1096GAT(408)
g369 and 1026GAT(394) 925GAT(332) ; 1108GAT(409)
g370 and 1031GAT(392) 925GAT(332) ; 1120GAT(410)
g371 and 996GAT(389) 873GAT(333) ; 1045GAT(411)
g372 and 1001GAT(387) 873GAT(333) ; 1057GAT(412)
g373 and 1006GAT(390) 873GAT(333) ; 1069GAT(413)
g374 and 1011GAT(388) 873GAT(333) ; 1081GAT(414)
g375 and 996GAT(389) 860GAT(334) ; 1042GAT(415)
g376 and 1001GAT(387) 860GAT(334) ; 1054GAT(416)
g377 and 1006GAT(390) 860GAT(334) ; 1066GAT(417)
g378 and 1011GAT(388) 860GAT(334) ; 1078GAT(418)
g379 and 996GAT(389) 847GAT(335) ; 1039GAT(419)
g380 and 1001GAT(387) 847GAT(335) ; 1051GAT(420)
g381 and 1006GAT(390) 847GAT(335) ; 1063GAT(421)
g382 and 1011GAT(388) 847GAT(335) ; 1075GAT(422)
g383 and 996GAT(389) 834GAT(336) ; 1036GAT(423)
g384 and 1001GAT(387) 834GAT(336) ; 1048GAT(424)
g385 and 1006GAT(390) 834GAT(336) ; 1060GAT(425)
g386 and 1011GAT(388) 834GAT(336) ; 1072GAT(426)
g387 and 1129GAT(398) 218GAT(31) ; 1225GAT(427)
g388 and 1126GAT(402) 211GAT(30) ; 1222GAT(428)
g389 and 1123GAT(406) 204GAT(29) ; 1219GAT(429)
g390 and 1120GAT(410) 197GAT(28) ; 1216GAT(430)
g391 and 1117GAT(397) 190GAT(27) ; 1213GAT(431)
g392 and 1114GAT(401) 183GAT(26) ; 1210GAT(432)
g393 and 1111GAT(405) 176GAT(25) ; 1207GAT(433)
g394 and 1108GAT(409) 169GAT(24) ; 1204GAT(434)
g395 and 1105GAT(396) 162GAT(23) ; 1201GAT(435)
g396 and 1102GAT(400) 155GAT(22) ; 1198GAT(436)
g397 and 1099GAT(404) 148GAT(21) ; 1195GAT(437)
g398 and 1096GAT(408) 141GAT(20) ; 1192GAT(438)
g399 and 1093GAT(395) 134GAT(19) ; 1189GAT(439)
g400 and 1090GAT(399) 127GAT(18) ; 1186GAT(440)
g401 and 1087GAT(403) 120GAT(17) ; 1183GAT(441)
g402 and 1084GAT(407) 113GAT(16) ; 1180GAT(442)
g403 and 1081GAT(414) 106GAT(15) ; 1177GAT(443)
g404 and 1078GAT(418) 99GAT(14) ; 1174GAT(444)
g405 and 1075GAT(422) 92GAT(13) ; 1171GAT(445)
g406 and 1072GAT(426) 85GAT(12) ; 1168GAT(446)
g407 and 1069GAT(413) 78GAT(11) ; 1165GAT(447)
g408 and 1066GAT(417) 71GAT(10) ; 1162GAT(448)
g409 and 1063GAT(421) 64GAT(9) ; 1159GAT(449)
g410 and 1060GAT(425) 57GAT(8) ; 1156GAT(450)
g411 and 1057GAT(412) 50GAT(7) ; 1153GAT(451)
g412 and 1054GAT(416) 43GAT(6) ; 1150GAT(452)
g413 and 1051GAT(420) 36GAT(5) ; 1147GAT(453)
g414 and 1048GAT(424) 29GAT(4) ; 1144GAT(454)
g415 and 1045GAT(411) 22GAT(3) ; 1141GAT(455)
g416 and 1042GAT(415) 15GAT(2) ; 1138GAT(456)
g417 and 1039GAT(419) 8GAT(1) ; 1135GAT(457)
g418 and 1036GAT(423) 1GAT(0) ; 1132GAT(458)
g419 and 1189GAT(439) 1093GAT(395) ; 1267GAT(459)
g420 and 1201GAT(435) 1105GAT(396) ; 1275GAT(460)
g421 and 1213GAT(431) 1117GAT(397) ; 1283GAT(461)
g422 and 1225GAT(427) 1129GAT(398) ; 1291GAT(462)
g423 and 1186GAT(440) 1090GAT(399) ; 1265GAT(463)
g424 and 1198GAT(436) 1102GAT(400) ; 1273GAT(464)
g425 and 1210GAT(432) 1114GAT(401) ; 1281GAT(465)
g426 and 1222GAT(428) 1126GAT(402) ; 1289GAT(466)
g427 and 1183GAT(441) 1087GAT(403) ; 1263GAT(467)
g428 and 1195GAT(437) 1099GAT(404) ; 1271GAT(468)
g429 and 1207GAT(433) 1111GAT(405) ; 1279GAT(469)
g430 and 1219GAT(429) 1123GAT(406) ; 1287GAT(470)
g431 and 1180GAT(442) 1084GAT(407) ; 1261GAT(471)
g432 and 1192GAT(438) 1096GAT(408) ; 1269GAT(472)
g433 and 1204GAT(434) 1108GAT(409) ; 1277GAT(473)
g434 and 1216GAT(430) 1120GAT(410) ; 1285GAT(474)
g435 and 1141GAT(455) 1045GAT(411) ; 1235GAT(475)
g436 and 1153GAT(451) 1057GAT(412) ; 1243GAT(476)
g437 and 1165GAT(447) 1069GAT(413) ; 1251GAT(477)
g438 and 1177GAT(443) 1081GAT(414) ; 1259GAT(478)
g439 and 1138GAT(456) 1042GAT(415) ; 1233GAT(479)
g440 and 1150GAT(452) 1054GAT(416) ; 1241GAT(480)
g441 and 1162GAT(448) 1066GAT(417) ; 1249GAT(481)
g442 and 1174GAT(444) 1078GAT(418) ; 1257GAT(482)
g443 and 1135GAT(457) 1039GAT(419) ; 1231GAT(483)
g444 and 1147GAT(453) 1051GAT(420) ; 1239GAT(484)
g445 and 1159GAT(449) 1063GAT(421) ; 1247GAT(485)
g446 and 1171GAT(445) 1075GAT(422) ; 1255GAT(486)
g447 and 1132GAT(458) 1036GAT(423) ; 1229GAT(487)
g448 and 1144GAT(454) 1048GAT(424) ; 1237GAT(488)
g449 and 1156GAT(450) 1060GAT(425) ; 1245GAT(489)
g450 and 1168GAT(446) 1072GAT(426) ; 1253GAT(490)
g451 and 1225GAT(427) 218GAT(31) ; 1290GAT(491)
g452 and 1222GAT(428) 211GAT(30) ; 1288GAT(492)
g453 and 1219GAT(429) 204GAT(29) ; 1286GAT(493)
g454 and 1216GAT(430) 197GAT(28) ; 1284GAT(494)
g455 and 1213GAT(431) 190GAT(27) ; 1282GAT(495)
g456 and 1210GAT(432) 183GAT(26) ; 1280GAT(496)
g457 and 1207GAT(433) 176GAT(25) ; 1278GAT(497)
g458 and 1204GAT(434) 169GAT(24) ; 1276GAT(498)
g459 and 1201GAT(435) 162GAT(23) ; 1274GAT(499)
g460 and 1198GAT(436) 155GAT(22) ; 1272GAT(500)
g461 and 1195GAT(437) 148GAT(21) ; 1270GAT(501)
g462 and 1192GAT(438) 141GAT(20) ; 1268GAT(502)
g463 and 1189GAT(439) 134GAT(19) ; 1266GAT(503)
g464 and 1186GAT(440) 127GAT(18) ; 1264GAT(504)
g465 and 1183GAT(441) 120GAT(17) ; 1262GAT(505)
g466 and 1180GAT(442) 113GAT(16) ; 1260GAT(506)
g467 and 1177GAT(443) 106GAT(15) ; 1258GAT(507)
g468 and 1174GAT(444) 99GAT(14) ; 1256GAT(508)
g469 and 1171GAT(445) 92GAT(13) ; 1254GAT(509)
g470 and 1168GAT(446) 85GAT(12) ; 1252GAT(510)
g471 and 1165GAT(447) 78GAT(11) ; 1250GAT(511)
g472 and 1162GAT(448) 71GAT(10) ; 1248GAT(512)
g473 and 1159GAT(449) 64GAT(9) ; 1246GAT(513)
g474 and 1156GAT(450) 57GAT(8) ; 1244GAT(514)
g475 and 1153GAT(451) 50GAT(7) ; 1242GAT(515)
g476 and 1150GAT(452) 43GAT(6) ; 1240GAT(516)
g477 and 1147GAT(453) 36GAT(5) ; 1238GAT(517)
g478 and 1144GAT(454) 29GAT(4) ; 1236GAT(518)
g479 and 1141GAT(455) 22GAT(3) ; 1234GAT(519)
g480 and 1138GAT(456) 15GAT(2) ; 1232GAT(520)
g481 and 1135GAT(457) 8GAT(1) ; 1230GAT(521)
g482 and 1132GAT(458) 1GAT(0) ; 1228GAT(522)
g483 and 1267GAT(459) 1266GAT(503) ; 1311GAT(523)
g484 and 1275GAT(460) 1274GAT(499) ; 1315GAT(524)
g485 and 1283GAT(461) 1282GAT(495) ; 1319GAT(525)
g486 and 1291GAT(462) 1290GAT(491) ; 1323GAT(526)
g487 and 1265GAT(463) 1264GAT(504) ; 1310GAT(527)
g488 and 1273GAT(464) 1272GAT(500) ; 1314GAT(528)
g489 and 1281GAT(465) 1280GAT(496) ; 1318GAT(529)
g490 and 1289GAT(466) 1288GAT(492) ; 1322GAT(530)
g491 and 1263GAT(467) 1262GAT(505) ; 1309GAT(531)
g492 and 1271GAT(468) 1270GAT(501) ; 1313GAT(532)
g493 and 1279GAT(469) 1278GAT(497) ; 1317GAT(533)
g494 and 1287GAT(470) 1286GAT(493) ; 1321GAT(534)
g495 and 1261GAT(471) 1260GAT(506) ; 1308GAT(535)
g496 and 1269GAT(472) 1268GAT(502) ; 1312GAT(536)
g497 and 1277GAT(473) 1276GAT(498) ; 1316GAT(537)
g498 and 1285GAT(474) 1284GAT(494) ; 1320GAT(538)
g499 and 1235GAT(475) 1234GAT(519) ; 1295GAT(539)
g500 and 1243GAT(476) 1242GAT(515) ; 1299GAT(540)
g501 and 1251GAT(477) 1250GAT(511) ; 1303GAT(541)
g502 and 1259GAT(478) 1258GAT(507) ; 1307GAT(542)
g503 and 1233GAT(479) 1232GAT(520) ; 1294GAT(543)
g504 and 1241GAT(480) 1240GAT(516) ; 1298GAT(544)
g505 and 1249GAT(481) 1248GAT(512) ; 1302GAT(545)
g506 and 1257GAT(482) 1256GAT(508) ; 1306GAT(546)
g507 and 1231GAT(483) 1230GAT(521) ; 1293GAT(547)
g508 and 1239GAT(484) 1238GAT(517) ; 1297GAT(548)
g509 and 1247GAT(485) 1246GAT(513) ; 1301GAT(549)
g510 and 1255GAT(486) 1254GAT(509) ; 1305GAT(550)
g511 and 1229GAT(487) 1228GAT(522) ; 1292GAT(551)
g512 and 1237GAT(488) 1236GAT(518) ; 1296GAT(552)
g513 and 1245GAT(489) 1244GAT(514) ; 1300GAT(553)
g514 and 1253GAT(490) 1252GAT(510) ; 1304GAT(554)
g515 and 1311GAT(523) ; 1343GAT(555)
g516 and 1315GAT(524) ; 1347GAT(556)
g517 and 1319GAT(525) ; 1351GAT(557)
g518 and 1323GAT(526) ; 1355GAT(558)
g519 and 1310GAT(527) ; 1342GAT(559)
g520 and 1314GAT(528) ; 1346GAT(560)
g521 and 1318GAT(529) ; 1350GAT(561)
g522 and 1322GAT(530) ; 1354GAT(562)
g523 and 1309GAT(531) ; 1341GAT(563)
g524 and 1313GAT(532) ; 1345GAT(564)
g525 and 1317GAT(533) ; 1349GAT(565)
g526 and 1321GAT(534) ; 1353GAT(566)
g527 and 1308GAT(535) ; 1340GAT(567)
g528 and 1312GAT(536) ; 1344GAT(568)
g529 and 1316GAT(537) ; 1348GAT(569)
g530 and 1320GAT(538) ; 1352GAT(570)
g531 and 1295GAT(539) ; 1327GAT(571)
g532 and 1299GAT(540) ; 1331GAT(572)
g533 and 1303GAT(541) ; 1335GAT(573)
g534 and 1307GAT(542) ; 1339GAT(574)
g535 and 1294GAT(543) ; 1326GAT(575)
g536 and 1298GAT(544) ; 1330GAT(576)
g537 and 1302GAT(545) ; 1334GAT(577)
g538 and 1306GAT(546) ; 1338GAT(578)
g539 and 1293GAT(547) ; 1325GAT(579)
g540 and 1297GAT(548) ; 1329GAT(580)
g541 and 1301GAT(549) ; 1333GAT(581)
g542 and 1305GAT(550) ; 1337GAT(582)
g543 and 1292GAT(551) ; 1324GAT(583)
g544 and 1296GAT(552) ; 1328GAT(584)
g545 and 1300GAT(553) ; 1332GAT(585)
g546 and 1304GAT(554) ; 1336GAT(586)
g547 not 982GAT(377) ; 982GAT(377)*
g548 not 983GAT(378) ; 983GAT(378)*
g549 not 984GAT(379) ; 984GAT(379)*
g550 not 985GAT(380) ; 985GAT(380)*
g551 not 978GAT(381) ; 978GAT(381)*
g552 not 979GAT(382) ; 979GAT(382)*
g553 not 980GAT(383) ; 980GAT(383)*
g554 not 981GAT(384) ; 981GAT(384)*
